magic
tech sky130A
magscale 1 2
timestamp 1715010268
<< nwell >>
rect -683 -584 683 584
<< pmos >>
rect -487 -436 -287 364
rect -229 -436 -29 364
rect 29 -436 229 364
rect 287 -436 487 364
<< pdiff >>
rect -545 321 -487 364
rect -545 287 -533 321
rect -499 287 -487 321
rect -545 253 -487 287
rect -545 219 -533 253
rect -499 219 -487 253
rect -545 185 -487 219
rect -545 151 -533 185
rect -499 151 -487 185
rect -545 117 -487 151
rect -545 83 -533 117
rect -499 83 -487 117
rect -545 49 -487 83
rect -545 15 -533 49
rect -499 15 -487 49
rect -545 -19 -487 15
rect -545 -53 -533 -19
rect -499 -53 -487 -19
rect -545 -87 -487 -53
rect -545 -121 -533 -87
rect -499 -121 -487 -87
rect -545 -155 -487 -121
rect -545 -189 -533 -155
rect -499 -189 -487 -155
rect -545 -223 -487 -189
rect -545 -257 -533 -223
rect -499 -257 -487 -223
rect -545 -291 -487 -257
rect -545 -325 -533 -291
rect -499 -325 -487 -291
rect -545 -359 -487 -325
rect -545 -393 -533 -359
rect -499 -393 -487 -359
rect -545 -436 -487 -393
rect -287 321 -229 364
rect -287 287 -275 321
rect -241 287 -229 321
rect -287 253 -229 287
rect -287 219 -275 253
rect -241 219 -229 253
rect -287 185 -229 219
rect -287 151 -275 185
rect -241 151 -229 185
rect -287 117 -229 151
rect -287 83 -275 117
rect -241 83 -229 117
rect -287 49 -229 83
rect -287 15 -275 49
rect -241 15 -229 49
rect -287 -19 -229 15
rect -287 -53 -275 -19
rect -241 -53 -229 -19
rect -287 -87 -229 -53
rect -287 -121 -275 -87
rect -241 -121 -229 -87
rect -287 -155 -229 -121
rect -287 -189 -275 -155
rect -241 -189 -229 -155
rect -287 -223 -229 -189
rect -287 -257 -275 -223
rect -241 -257 -229 -223
rect -287 -291 -229 -257
rect -287 -325 -275 -291
rect -241 -325 -229 -291
rect -287 -359 -229 -325
rect -287 -393 -275 -359
rect -241 -393 -229 -359
rect -287 -436 -229 -393
rect -29 321 29 364
rect -29 287 -17 321
rect 17 287 29 321
rect -29 253 29 287
rect -29 219 -17 253
rect 17 219 29 253
rect -29 185 29 219
rect -29 151 -17 185
rect 17 151 29 185
rect -29 117 29 151
rect -29 83 -17 117
rect 17 83 29 117
rect -29 49 29 83
rect -29 15 -17 49
rect 17 15 29 49
rect -29 -19 29 15
rect -29 -53 -17 -19
rect 17 -53 29 -19
rect -29 -87 29 -53
rect -29 -121 -17 -87
rect 17 -121 29 -87
rect -29 -155 29 -121
rect -29 -189 -17 -155
rect 17 -189 29 -155
rect -29 -223 29 -189
rect -29 -257 -17 -223
rect 17 -257 29 -223
rect -29 -291 29 -257
rect -29 -325 -17 -291
rect 17 -325 29 -291
rect -29 -359 29 -325
rect -29 -393 -17 -359
rect 17 -393 29 -359
rect -29 -436 29 -393
rect 229 321 287 364
rect 229 287 241 321
rect 275 287 287 321
rect 229 253 287 287
rect 229 219 241 253
rect 275 219 287 253
rect 229 185 287 219
rect 229 151 241 185
rect 275 151 287 185
rect 229 117 287 151
rect 229 83 241 117
rect 275 83 287 117
rect 229 49 287 83
rect 229 15 241 49
rect 275 15 287 49
rect 229 -19 287 15
rect 229 -53 241 -19
rect 275 -53 287 -19
rect 229 -87 287 -53
rect 229 -121 241 -87
rect 275 -121 287 -87
rect 229 -155 287 -121
rect 229 -189 241 -155
rect 275 -189 287 -155
rect 229 -223 287 -189
rect 229 -257 241 -223
rect 275 -257 287 -223
rect 229 -291 287 -257
rect 229 -325 241 -291
rect 275 -325 287 -291
rect 229 -359 287 -325
rect 229 -393 241 -359
rect 275 -393 287 -359
rect 229 -436 287 -393
rect 487 321 545 364
rect 487 287 499 321
rect 533 287 545 321
rect 487 253 545 287
rect 487 219 499 253
rect 533 219 545 253
rect 487 185 545 219
rect 487 151 499 185
rect 533 151 545 185
rect 487 117 545 151
rect 487 83 499 117
rect 533 83 545 117
rect 487 49 545 83
rect 487 15 499 49
rect 533 15 545 49
rect 487 -19 545 15
rect 487 -53 499 -19
rect 533 -53 545 -19
rect 487 -87 545 -53
rect 487 -121 499 -87
rect 533 -121 545 -87
rect 487 -155 545 -121
rect 487 -189 499 -155
rect 533 -189 545 -155
rect 487 -223 545 -189
rect 487 -257 499 -223
rect 533 -257 545 -223
rect 487 -291 545 -257
rect 487 -325 499 -291
rect 533 -325 545 -291
rect 487 -359 545 -325
rect 487 -393 499 -359
rect 533 -393 545 -359
rect 487 -436 545 -393
<< pdiffc >>
rect -533 287 -499 321
rect -533 219 -499 253
rect -533 151 -499 185
rect -533 83 -499 117
rect -533 15 -499 49
rect -533 -53 -499 -19
rect -533 -121 -499 -87
rect -533 -189 -499 -155
rect -533 -257 -499 -223
rect -533 -325 -499 -291
rect -533 -393 -499 -359
rect -275 287 -241 321
rect -275 219 -241 253
rect -275 151 -241 185
rect -275 83 -241 117
rect -275 15 -241 49
rect -275 -53 -241 -19
rect -275 -121 -241 -87
rect -275 -189 -241 -155
rect -275 -257 -241 -223
rect -275 -325 -241 -291
rect -275 -393 -241 -359
rect -17 287 17 321
rect -17 219 17 253
rect -17 151 17 185
rect -17 83 17 117
rect -17 15 17 49
rect -17 -53 17 -19
rect -17 -121 17 -87
rect -17 -189 17 -155
rect -17 -257 17 -223
rect -17 -325 17 -291
rect -17 -393 17 -359
rect 241 287 275 321
rect 241 219 275 253
rect 241 151 275 185
rect 241 83 275 117
rect 241 15 275 49
rect 241 -53 275 -19
rect 241 -121 275 -87
rect 241 -189 275 -155
rect 241 -257 275 -223
rect 241 -325 275 -291
rect 241 -393 275 -359
rect 499 287 533 321
rect 499 219 533 253
rect 499 151 533 185
rect 499 83 533 117
rect 499 15 533 49
rect 499 -53 533 -19
rect 499 -121 533 -87
rect 499 -189 533 -155
rect 499 -257 533 -223
rect 499 -325 533 -291
rect 499 -393 533 -359
<< nsubdiff >>
rect -647 514 -527 548
rect -493 514 -459 548
rect -425 514 -391 548
rect -357 514 -323 548
rect -289 514 -255 548
rect -221 514 -187 548
rect -153 514 -119 548
rect -85 514 -51 548
rect -17 514 17 548
rect 51 514 85 548
rect 119 514 153 548
rect 187 514 221 548
rect 255 514 289 548
rect 323 514 357 548
rect 391 514 425 548
rect 459 514 493 548
rect 527 514 647 548
rect -647 425 -613 514
rect -647 357 -613 391
rect 613 425 647 514
rect -647 289 -613 323
rect -647 221 -613 255
rect -647 153 -613 187
rect -647 85 -613 119
rect -647 17 -613 51
rect -647 -51 -613 -17
rect -647 -119 -613 -85
rect -647 -187 -613 -153
rect -647 -255 -613 -221
rect -647 -323 -613 -289
rect -647 -391 -613 -357
rect -647 -514 -613 -425
rect 613 357 647 391
rect 613 289 647 323
rect 613 221 647 255
rect 613 153 647 187
rect 613 85 647 119
rect 613 17 647 51
rect 613 -51 647 -17
rect 613 -119 647 -85
rect 613 -187 647 -153
rect 613 -255 647 -221
rect 613 -323 647 -289
rect 613 -391 647 -357
rect 613 -514 647 -425
rect -647 -548 -527 -514
rect -493 -548 -459 -514
rect -425 -548 -391 -514
rect -357 -548 -323 -514
rect -289 -548 -255 -514
rect -221 -548 -187 -514
rect -153 -548 -119 -514
rect -85 -548 -51 -514
rect -17 -548 17 -514
rect 51 -548 85 -514
rect 119 -548 153 -514
rect 187 -548 221 -514
rect 255 -548 289 -514
rect 323 -548 357 -514
rect 391 -548 425 -514
rect 459 -548 493 -514
rect 527 -548 647 -514
<< nsubdiffcont >>
rect -527 514 -493 548
rect -459 514 -425 548
rect -391 514 -357 548
rect -323 514 -289 548
rect -255 514 -221 548
rect -187 514 -153 548
rect -119 514 -85 548
rect -51 514 -17 548
rect 17 514 51 548
rect 85 514 119 548
rect 153 514 187 548
rect 221 514 255 548
rect 289 514 323 548
rect 357 514 391 548
rect 425 514 459 548
rect 493 514 527 548
rect -647 391 -613 425
rect 613 391 647 425
rect -647 323 -613 357
rect -647 255 -613 289
rect -647 187 -613 221
rect -647 119 -613 153
rect -647 51 -613 85
rect -647 -17 -613 17
rect -647 -85 -613 -51
rect -647 -153 -613 -119
rect -647 -221 -613 -187
rect -647 -289 -613 -255
rect -647 -357 -613 -323
rect -647 -425 -613 -391
rect 613 323 647 357
rect 613 255 647 289
rect 613 187 647 221
rect 613 119 647 153
rect 613 51 647 85
rect 613 -17 647 17
rect 613 -85 647 -51
rect 613 -153 647 -119
rect 613 -221 647 -187
rect 613 -289 647 -255
rect 613 -357 647 -323
rect 613 -425 647 -391
rect -527 -548 -493 -514
rect -459 -548 -425 -514
rect -391 -548 -357 -514
rect -323 -548 -289 -514
rect -255 -548 -221 -514
rect -187 -548 -153 -514
rect -119 -548 -85 -514
rect -51 -548 -17 -514
rect 17 -548 51 -514
rect 85 -548 119 -514
rect 153 -548 187 -514
rect 221 -548 255 -514
rect 289 -548 323 -514
rect 357 -548 391 -514
rect 425 -548 459 -514
rect 493 -548 527 -514
<< poly >>
rect -487 445 -287 461
rect -487 411 -438 445
rect -404 411 -370 445
rect -336 411 -287 445
rect -487 364 -287 411
rect -229 445 -29 461
rect -229 411 -180 445
rect -146 411 -112 445
rect -78 411 -29 445
rect -229 364 -29 411
rect 29 445 229 461
rect 29 411 78 445
rect 112 411 146 445
rect 180 411 229 445
rect 29 364 229 411
rect 287 445 487 461
rect 287 411 336 445
rect 370 411 404 445
rect 438 411 487 445
rect 287 364 487 411
rect -487 -462 -287 -436
rect -229 -462 -29 -436
rect 29 -462 229 -436
rect 287 -462 487 -436
<< polycont >>
rect -438 411 -404 445
rect -370 411 -336 445
rect -180 411 -146 445
rect -112 411 -78 445
rect 78 411 112 445
rect 146 411 180 445
rect 336 411 370 445
rect 404 411 438 445
<< locali >>
rect -647 514 -527 548
rect -493 514 -459 548
rect -425 514 -391 548
rect -357 514 -323 548
rect -289 514 -255 548
rect -221 514 -187 548
rect -153 514 -119 548
rect -85 514 -51 548
rect -17 514 17 548
rect 51 514 85 548
rect 119 514 153 548
rect 187 514 221 548
rect 255 514 289 548
rect 323 514 357 548
rect 391 514 425 548
rect 459 514 493 548
rect 527 514 647 548
rect -647 425 -613 514
rect -487 411 -440 445
rect -404 411 -370 445
rect -334 411 -287 445
rect -229 411 -182 445
rect -146 411 -112 445
rect -76 411 -29 445
rect 29 411 76 445
rect 112 411 146 445
rect 182 411 229 445
rect 287 411 334 445
rect 370 411 404 445
rect 440 411 487 445
rect 613 425 647 514
rect -647 357 -613 391
rect -647 289 -613 323
rect -647 221 -613 255
rect -647 153 -613 187
rect -647 85 -613 119
rect -647 17 -613 51
rect -647 -51 -613 -17
rect -647 -119 -613 -85
rect -647 -187 -613 -153
rect -647 -255 -613 -221
rect -647 -323 -613 -289
rect -647 -391 -613 -357
rect -647 -514 -613 -425
rect -533 341 -499 368
rect -533 269 -499 287
rect -533 197 -499 219
rect -533 125 -499 151
rect -533 53 -499 83
rect -533 -19 -499 15
rect -533 -87 -499 -53
rect -533 -155 -499 -125
rect -533 -223 -499 -197
rect -533 -291 -499 -269
rect -533 -359 -499 -341
rect -533 -440 -499 -413
rect -275 341 -241 368
rect -275 269 -241 287
rect -275 197 -241 219
rect -275 125 -241 151
rect -275 53 -241 83
rect -275 -19 -241 15
rect -275 -87 -241 -53
rect -275 -155 -241 -125
rect -275 -223 -241 -197
rect -275 -291 -241 -269
rect -275 -359 -241 -341
rect -275 -440 -241 -413
rect -17 341 17 368
rect -17 269 17 287
rect -17 197 17 219
rect -17 125 17 151
rect -17 53 17 83
rect -17 -19 17 15
rect -17 -87 17 -53
rect -17 -155 17 -125
rect -17 -223 17 -197
rect -17 -291 17 -269
rect -17 -359 17 -341
rect -17 -440 17 -413
rect 241 341 275 368
rect 241 269 275 287
rect 241 197 275 219
rect 241 125 275 151
rect 241 53 275 83
rect 241 -19 275 15
rect 241 -87 275 -53
rect 241 -155 275 -125
rect 241 -223 275 -197
rect 241 -291 275 -269
rect 241 -359 275 -341
rect 241 -440 275 -413
rect 499 341 533 368
rect 499 269 533 287
rect 499 197 533 219
rect 499 125 533 151
rect 499 53 533 83
rect 499 -19 533 15
rect 499 -87 533 -53
rect 499 -155 533 -125
rect 499 -223 533 -197
rect 499 -291 533 -269
rect 499 -359 533 -341
rect 499 -440 533 -413
rect 613 357 647 391
rect 613 289 647 323
rect 613 221 647 255
rect 613 153 647 187
rect 613 85 647 119
rect 613 17 647 51
rect 613 -51 647 -17
rect 613 -119 647 -85
rect 613 -187 647 -153
rect 613 -255 647 -221
rect 613 -323 647 -289
rect 613 -391 647 -357
rect 613 -514 647 -425
rect -647 -548 -527 -514
rect -493 -548 -459 -514
rect -425 -548 -391 -514
rect -357 -548 -323 -514
rect -289 -548 -255 -514
rect -221 -548 -187 -514
rect -153 -548 -119 -514
rect -85 -548 -51 -514
rect -17 -548 17 -514
rect 51 -548 85 -514
rect 119 -548 153 -514
rect 187 -548 221 -514
rect 255 -548 289 -514
rect 323 -548 357 -514
rect 391 -548 425 -514
rect 459 -548 493 -514
rect 527 -548 647 -514
<< viali >>
rect -440 411 -438 445
rect -438 411 -406 445
rect -368 411 -336 445
rect -336 411 -334 445
rect -182 411 -180 445
rect -180 411 -148 445
rect -110 411 -78 445
rect -78 411 -76 445
rect 76 411 78 445
rect 78 411 110 445
rect 148 411 180 445
rect 180 411 182 445
rect 334 411 336 445
rect 336 411 368 445
rect 406 411 438 445
rect 438 411 440 445
rect -533 321 -499 341
rect -533 307 -499 321
rect -533 253 -499 269
rect -533 235 -499 253
rect -533 185 -499 197
rect -533 163 -499 185
rect -533 117 -499 125
rect -533 91 -499 117
rect -533 49 -499 53
rect -533 19 -499 49
rect -533 -53 -499 -19
rect -533 -121 -499 -91
rect -533 -125 -499 -121
rect -533 -189 -499 -163
rect -533 -197 -499 -189
rect -533 -257 -499 -235
rect -533 -269 -499 -257
rect -533 -325 -499 -307
rect -533 -341 -499 -325
rect -533 -393 -499 -379
rect -533 -413 -499 -393
rect -275 321 -241 341
rect -275 307 -241 321
rect -275 253 -241 269
rect -275 235 -241 253
rect -275 185 -241 197
rect -275 163 -241 185
rect -275 117 -241 125
rect -275 91 -241 117
rect -275 49 -241 53
rect -275 19 -241 49
rect -275 -53 -241 -19
rect -275 -121 -241 -91
rect -275 -125 -241 -121
rect -275 -189 -241 -163
rect -275 -197 -241 -189
rect -275 -257 -241 -235
rect -275 -269 -241 -257
rect -275 -325 -241 -307
rect -275 -341 -241 -325
rect -275 -393 -241 -379
rect -275 -413 -241 -393
rect -17 321 17 341
rect -17 307 17 321
rect -17 253 17 269
rect -17 235 17 253
rect -17 185 17 197
rect -17 163 17 185
rect -17 117 17 125
rect -17 91 17 117
rect -17 49 17 53
rect -17 19 17 49
rect -17 -53 17 -19
rect -17 -121 17 -91
rect -17 -125 17 -121
rect -17 -189 17 -163
rect -17 -197 17 -189
rect -17 -257 17 -235
rect -17 -269 17 -257
rect -17 -325 17 -307
rect -17 -341 17 -325
rect -17 -393 17 -379
rect -17 -413 17 -393
rect 241 321 275 341
rect 241 307 275 321
rect 241 253 275 269
rect 241 235 275 253
rect 241 185 275 197
rect 241 163 275 185
rect 241 117 275 125
rect 241 91 275 117
rect 241 49 275 53
rect 241 19 275 49
rect 241 -53 275 -19
rect 241 -121 275 -91
rect 241 -125 275 -121
rect 241 -189 275 -163
rect 241 -197 275 -189
rect 241 -257 275 -235
rect 241 -269 275 -257
rect 241 -325 275 -307
rect 241 -341 275 -325
rect 241 -393 275 -379
rect 241 -413 275 -393
rect 499 321 533 341
rect 499 307 533 321
rect 499 253 533 269
rect 499 235 533 253
rect 499 185 533 197
rect 499 163 533 185
rect 499 117 533 125
rect 499 91 533 117
rect 499 49 533 53
rect 499 19 533 49
rect 499 -53 533 -19
rect 499 -121 533 -91
rect 499 -125 533 -121
rect 499 -189 533 -163
rect 499 -197 533 -189
rect 499 -257 533 -235
rect 499 -269 533 -257
rect 499 -325 533 -307
rect 499 -341 533 -325
rect 499 -393 533 -379
rect 499 -413 533 -393
<< metal1 >>
rect -483 445 -291 451
rect -483 411 -440 445
rect -406 411 -368 445
rect -334 411 -291 445
rect -483 405 -291 411
rect -225 445 -33 451
rect -225 411 -182 445
rect -148 411 -110 445
rect -76 411 -33 445
rect -225 405 -33 411
rect 33 445 225 451
rect 33 411 76 445
rect 110 411 148 445
rect 182 411 225 445
rect 33 405 225 411
rect 291 445 483 451
rect 291 411 334 445
rect 368 411 406 445
rect 440 411 483 445
rect 291 405 483 411
rect -539 341 -493 364
rect -539 307 -533 341
rect -499 307 -493 341
rect -539 269 -493 307
rect -539 235 -533 269
rect -499 235 -493 269
rect -539 197 -493 235
rect -539 163 -533 197
rect -499 163 -493 197
rect -539 125 -493 163
rect -539 91 -533 125
rect -499 91 -493 125
rect -539 53 -493 91
rect -539 19 -533 53
rect -499 19 -493 53
rect -539 -19 -493 19
rect -539 -53 -533 -19
rect -499 -53 -493 -19
rect -539 -91 -493 -53
rect -539 -125 -533 -91
rect -499 -125 -493 -91
rect -539 -163 -493 -125
rect -539 -197 -533 -163
rect -499 -197 -493 -163
rect -539 -235 -493 -197
rect -539 -269 -533 -235
rect -499 -269 -493 -235
rect -539 -307 -493 -269
rect -539 -341 -533 -307
rect -499 -341 -493 -307
rect -539 -379 -493 -341
rect -539 -413 -533 -379
rect -499 -413 -493 -379
rect -539 -436 -493 -413
rect -281 341 -235 364
rect -281 307 -275 341
rect -241 307 -235 341
rect -281 269 -235 307
rect -281 235 -275 269
rect -241 235 -235 269
rect -281 197 -235 235
rect -281 163 -275 197
rect -241 163 -235 197
rect -281 125 -235 163
rect -281 91 -275 125
rect -241 91 -235 125
rect -281 53 -235 91
rect -281 19 -275 53
rect -241 19 -235 53
rect -281 -19 -235 19
rect -281 -53 -275 -19
rect -241 -53 -235 -19
rect -281 -91 -235 -53
rect -281 -125 -275 -91
rect -241 -125 -235 -91
rect -281 -163 -235 -125
rect -281 -197 -275 -163
rect -241 -197 -235 -163
rect -281 -235 -235 -197
rect -281 -269 -275 -235
rect -241 -269 -235 -235
rect -281 -307 -235 -269
rect -281 -341 -275 -307
rect -241 -341 -235 -307
rect -281 -379 -235 -341
rect -281 -413 -275 -379
rect -241 -413 -235 -379
rect -281 -436 -235 -413
rect -23 341 23 364
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -436 23 -413
rect 235 341 281 364
rect 235 307 241 341
rect 275 307 281 341
rect 235 269 281 307
rect 235 235 241 269
rect 275 235 281 269
rect 235 197 281 235
rect 235 163 241 197
rect 275 163 281 197
rect 235 125 281 163
rect 235 91 241 125
rect 275 91 281 125
rect 235 53 281 91
rect 235 19 241 53
rect 275 19 281 53
rect 235 -19 281 19
rect 235 -53 241 -19
rect 275 -53 281 -19
rect 235 -91 281 -53
rect 235 -125 241 -91
rect 275 -125 281 -91
rect 235 -163 281 -125
rect 235 -197 241 -163
rect 275 -197 281 -163
rect 235 -235 281 -197
rect 235 -269 241 -235
rect 275 -269 281 -235
rect 235 -307 281 -269
rect 235 -341 241 -307
rect 275 -341 281 -307
rect 235 -379 281 -341
rect 235 -413 241 -379
rect 275 -413 281 -379
rect 235 -436 281 -413
rect 493 341 539 364
rect 493 307 499 341
rect 533 307 539 341
rect 493 269 539 307
rect 493 235 499 269
rect 533 235 539 269
rect 493 197 539 235
rect 493 163 499 197
rect 533 163 539 197
rect 493 125 539 163
rect 493 91 499 125
rect 533 91 539 125
rect 493 53 539 91
rect 493 19 499 53
rect 533 19 539 53
rect 493 -19 539 19
rect 493 -53 499 -19
rect 533 -53 539 -19
rect 493 -91 539 -53
rect 493 -125 499 -91
rect 533 -125 539 -91
rect 493 -163 539 -125
rect 493 -197 499 -163
rect 533 -197 539 -163
rect 493 -235 539 -197
rect 493 -269 499 -235
rect 533 -269 539 -235
rect 493 -307 539 -269
rect 493 -341 499 -307
rect 533 -341 539 -307
rect 493 -379 539 -341
rect 493 -413 499 -379
rect 533 -413 539 -379
rect 493 -436 539 -413
<< properties >>
string FIXED_BBOX -630 -531 630 531
<< end >>
