magic
tech sky130A
magscale 1 2
timestamp 1715625863
<< error_p >>
rect -458 -131 -400 69
rect 400 -131 458 69
<< pwell >>
rect -484 -157 484 95
<< nmoslvt >>
rect -400 -131 400 69
<< ndiff >>
rect -458 54 -400 69
rect -458 20 -446 54
rect -412 20 -400 54
rect -458 -14 -400 20
rect -458 -48 -446 -14
rect -412 -48 -400 -14
rect -458 -82 -400 -48
rect -458 -116 -446 -82
rect -412 -116 -400 -82
rect -458 -131 -400 -116
rect 400 54 458 69
rect 400 20 412 54
rect 446 20 458 54
rect 400 -14 458 20
rect 400 -48 412 -14
rect 446 -48 458 -14
rect 400 -82 458 -48
rect 400 -116 412 -82
rect 446 -116 458 -82
rect 400 -131 458 -116
<< ndiffc >>
rect -446 20 -412 54
rect -446 -48 -412 -14
rect -446 -116 -412 -82
rect 412 20 446 54
rect 412 -48 446 -14
rect 412 -116 446 -82
<< poly >>
rect -400 141 400 157
rect -400 107 -357 141
rect -323 107 -289 141
rect -255 107 -221 141
rect -187 107 -153 141
rect -119 107 -85 141
rect -51 107 -17 141
rect 17 107 51 141
rect 85 107 119 141
rect 153 107 187 141
rect 221 107 255 141
rect 289 107 323 141
rect 357 107 400 141
rect -400 69 400 107
rect -400 -157 400 -131
<< polycont >>
rect -357 107 -323 141
rect -289 107 -255 141
rect -221 107 -187 141
rect -153 107 -119 141
rect -85 107 -51 141
rect -17 107 17 141
rect 51 107 85 141
rect 119 107 153 141
rect 187 107 221 141
rect 255 107 289 141
rect 323 107 357 141
<< locali >>
rect -400 107 -377 141
rect -323 107 -305 141
rect -255 107 -233 141
rect -187 107 -161 141
rect -119 107 -89 141
rect -51 107 -17 141
rect 17 107 51 141
rect 89 107 119 141
rect 161 107 187 141
rect 233 107 255 141
rect 305 107 323 141
rect 377 107 400 141
rect -446 54 -412 73
rect -446 -14 -412 -12
rect -446 -50 -412 -48
rect -446 -135 -412 -116
rect 412 54 446 73
rect 412 -14 446 -12
rect 412 -50 446 -48
rect 412 -135 446 -116
<< viali >>
rect -377 107 -357 141
rect -357 107 -343 141
rect -305 107 -289 141
rect -289 107 -271 141
rect -233 107 -221 141
rect -221 107 -199 141
rect -161 107 -153 141
rect -153 107 -127 141
rect -89 107 -85 141
rect -85 107 -55 141
rect -17 107 17 141
rect 55 107 85 141
rect 85 107 89 141
rect 127 107 153 141
rect 153 107 161 141
rect 199 107 221 141
rect 221 107 233 141
rect 271 107 289 141
rect 289 107 305 141
rect 343 107 357 141
rect 357 107 377 141
rect -446 20 -412 22
rect -446 -12 -412 20
rect -446 -82 -412 -50
rect -446 -84 -412 -82
rect 412 20 446 22
rect 412 -12 446 20
rect 412 -82 446 -50
rect 412 -84 446 -82
<< metal1 >>
rect -396 141 396 147
rect -396 107 -377 141
rect -343 107 -305 141
rect -271 107 -233 141
rect -199 107 -161 141
rect -127 107 -89 141
rect -55 107 -17 141
rect 17 107 55 141
rect 89 107 127 141
rect 161 107 199 141
rect 233 107 271 141
rect 305 107 343 141
rect 377 107 396 141
rect -396 101 396 107
rect -452 22 -406 69
rect -452 -12 -446 22
rect -412 -12 -406 22
rect -452 -50 -406 -12
rect -452 -84 -446 -50
rect -412 -84 -406 -50
rect -452 -131 -406 -84
rect 406 22 452 69
rect 406 -12 412 22
rect 446 -12 452 22
rect 406 -50 452 -12
rect 406 -84 412 -50
rect 446 -84 452 -50
rect 406 -131 452 -84
<< end >>
