magic
tech sky130A
magscale 1 2
timestamp 1715616696
<< pwell >>
rect -274 -1462 270 1364
<< psubdiff >>
rect -86 -1459 114 -1425
<< xpolycontact >>
rect -194 846 -124 1282
rect -194 -1282 -124 -846
rect 124 846 194 1282
rect 124 -1282 194 -846
<< xpolyres >>
rect -194 -846 -124 846
rect 124 -846 194 846
<< viali >>
rect -176 1228 -142 1262
rect -176 1156 -142 1190
rect -176 1084 -142 1118
rect -176 1012 -142 1046
rect -176 940 -142 974
rect -176 868 -142 902
rect 142 1228 176 1262
rect 142 1156 176 1190
rect 142 1084 176 1118
rect 142 1012 176 1046
rect 142 940 176 974
rect 142 868 176 902
rect -176 -903 -142 -869
rect -176 -975 -142 -941
rect -176 -1047 -142 -1013
rect -176 -1119 -142 -1085
rect -176 -1191 -142 -1157
rect -176 -1263 -142 -1229
rect 142 -903 176 -869
rect 142 -975 176 -941
rect 142 -1047 176 -1013
rect 142 -1119 176 -1085
rect 142 -1191 176 -1157
rect 142 -1263 176 -1229
<< metal1 >>
rect -184 1262 -134 1276
rect -184 1228 -176 1262
rect -142 1228 -134 1262
rect -184 1190 -134 1228
rect -184 1156 -176 1190
rect -142 1156 -134 1190
rect -184 1118 -134 1156
rect -184 1084 -176 1118
rect -142 1084 -134 1118
rect -184 1046 -134 1084
rect -184 1012 -176 1046
rect -142 1012 -134 1046
rect -184 974 -134 1012
rect -184 940 -176 974
rect -142 940 -134 974
rect -184 902 -134 940
rect -184 868 -176 902
rect -142 868 -134 902
rect -184 855 -134 868
rect 134 1262 184 1276
rect 134 1228 142 1262
rect 176 1228 184 1262
rect 134 1190 184 1228
rect 134 1156 142 1190
rect 176 1156 184 1190
rect 134 1118 184 1156
rect 134 1084 142 1118
rect 176 1084 184 1118
rect 134 1046 184 1084
rect 134 1012 142 1046
rect 176 1012 184 1046
rect 134 974 184 1012
rect 134 940 142 974
rect 176 940 184 974
rect 134 902 184 940
rect 134 868 142 902
rect 176 868 184 902
rect 134 855 184 868
rect -184 -869 -134 -855
rect -184 -903 -176 -869
rect -142 -903 -134 -869
rect -184 -941 -134 -903
rect -184 -975 -176 -941
rect -142 -975 -134 -941
rect -184 -1013 -134 -975
rect -184 -1047 -176 -1013
rect -142 -1047 -134 -1013
rect -184 -1085 -134 -1047
rect -184 -1119 -176 -1085
rect -142 -1119 -134 -1085
rect -184 -1157 -134 -1119
rect -184 -1191 -176 -1157
rect -142 -1191 -134 -1157
rect -184 -1229 -134 -1191
rect -184 -1263 -176 -1229
rect -142 -1263 -134 -1229
rect -184 -1276 -134 -1263
rect 134 -869 184 -855
rect 134 -903 142 -869
rect 176 -903 184 -869
rect 134 -941 184 -903
rect 134 -975 142 -941
rect 176 -975 184 -941
rect 134 -1013 184 -975
rect 134 -1047 142 -1013
rect 176 -1047 184 -1013
rect 134 -1085 184 -1047
rect 134 -1119 142 -1085
rect 176 -1119 184 -1085
rect 134 -1157 184 -1119
rect 134 -1191 142 -1157
rect 176 -1191 184 -1157
rect 134 -1229 184 -1191
rect 134 -1263 142 -1229
rect 176 -1263 184 -1229
rect 134 -1276 184 -1263
<< end >>
