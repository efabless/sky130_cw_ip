magic
tech sky130A
magscale 1 2
timestamp 1715010268
<< nwell >>
rect -194 -198 194 126
<< pmoslvt >>
rect -100 -136 100 64
<< pdiff >>
rect -158 49 -100 64
rect -158 15 -146 49
rect -112 15 -100 49
rect -158 -19 -100 15
rect -158 -53 -146 -19
rect -112 -53 -100 -19
rect -158 -87 -100 -53
rect -158 -121 -146 -87
rect -112 -121 -100 -87
rect -158 -136 -100 -121
rect 100 49 158 64
rect 100 15 112 49
rect 146 15 158 49
rect 100 -19 158 15
rect 100 -53 112 -19
rect 146 -53 158 -19
rect 100 -87 158 -53
rect 100 -121 112 -87
rect 146 -121 158 -87
rect 100 -136 158 -121
<< pdiffc >>
rect -146 15 -112 49
rect -146 -53 -112 -19
rect -146 -121 -112 -87
rect 112 15 146 49
rect 112 -53 146 -19
rect 112 -121 146 -87
<< poly >>
rect -100 64 100 90
rect -100 -162 100 -136
<< locali >>
rect -146 49 -112 68
rect -146 -19 -112 -17
rect -146 -55 -112 -53
rect -146 -140 -112 -121
rect 112 49 146 68
rect 112 -19 146 -17
rect 112 -55 146 -53
rect 112 -140 146 -121
<< viali >>
rect -146 15 -112 17
rect -146 -17 -112 15
rect -146 -87 -112 -55
rect -146 -89 -112 -87
rect 112 15 146 17
rect 112 -17 146 15
rect 112 -87 146 -55
rect 112 -89 146 -87
<< metal1 >>
rect -152 17 -106 64
rect -152 -17 -146 17
rect -112 -17 -106 17
rect -152 -55 -106 -17
rect -152 -89 -146 -55
rect -112 -89 -106 -55
rect -152 -136 -106 -89
rect 106 17 152 64
rect 106 -17 112 17
rect 146 -17 152 17
rect 106 -55 152 -17
rect 106 -89 112 -55
rect 146 -89 152 -55
rect 106 -136 152 -89
<< end >>
