magic
tech sky130A
magscale 1 2
timestamp 1715625863
<< nwell >>
rect -11408 12081 -8946 16692
<< nsubdiff >>
rect -11372 16622 -11285 16656
rect -11251 16622 -11217 16656
rect -11183 16622 -11149 16656
rect -11115 16622 -11081 16656
rect -11047 16622 -11013 16656
rect -10979 16622 -10945 16656
rect -10911 16622 -10877 16656
rect -10843 16622 -10809 16656
rect -10775 16622 -10741 16656
rect -10707 16622 -10673 16656
rect -10639 16622 -10605 16656
rect -10571 16622 -10537 16656
rect -10503 16622 -10469 16656
rect -10435 16622 -10401 16656
rect -10367 16622 -10333 16656
rect -10299 16622 -10265 16656
rect -10231 16622 -10197 16656
rect -10163 16622 -10129 16656
rect -10095 16622 -10061 16656
rect -10027 16622 -9993 16656
rect -9959 16622 -9925 16656
rect -9891 16622 -9857 16656
rect -9823 16622 -9789 16656
rect -9755 16622 -9721 16656
rect -9687 16622 -9653 16656
rect -9619 16622 -9585 16656
rect -9551 16622 -9517 16656
rect -9483 16622 -9449 16656
rect -9415 16622 -9381 16656
rect -9347 16622 -9313 16656
rect -9279 16622 -9245 16656
rect -9211 16622 -9177 16656
rect -9143 16622 -8982 16656
rect -11372 16516 -11338 16622
rect -11372 16448 -11338 16482
rect -11372 16380 -11338 16414
rect -11372 16312 -11338 16346
rect -11372 16244 -11338 16278
rect -11372 16176 -11338 16210
rect -11372 16108 -11338 16142
rect -11372 16040 -11338 16074
rect -11372 15972 -11338 16006
rect -11372 15904 -11338 15938
rect -11372 15836 -11338 15870
rect -11372 15768 -11338 15802
rect -11372 15700 -11338 15734
rect -11372 15632 -11338 15666
rect -11372 15564 -11338 15598
rect -11372 15496 -11338 15530
rect -11372 15428 -11338 15462
rect -11372 15360 -11338 15394
rect -11372 15292 -11338 15326
rect -11372 15224 -11338 15258
rect -11372 15156 -11338 15190
rect -11372 15088 -11338 15122
rect -11372 15020 -11338 15054
rect -11372 14952 -11338 14986
rect -11372 14884 -11338 14918
rect -11372 14816 -11338 14850
rect -11372 14748 -11338 14782
rect -11372 14680 -11338 14714
rect -11372 14612 -11338 14646
rect -11372 14544 -11338 14578
rect -11372 14476 -11338 14510
rect -11372 14408 -11338 14442
rect -11372 14340 -11338 14374
rect -11372 14272 -11338 14306
rect -11372 14204 -11338 14238
rect -11372 14136 -11338 14170
rect -11372 14068 -11338 14102
rect -11372 14000 -11338 14034
rect -11372 13932 -11338 13966
rect -11372 13864 -11338 13898
rect -11372 13796 -11338 13830
rect -11372 13728 -11338 13762
rect -11372 13660 -11338 13694
rect -11372 13592 -11338 13626
rect -11372 13524 -11338 13558
rect -11372 13456 -11338 13490
rect -11372 13388 -11338 13422
rect -11372 13320 -11338 13354
rect -11372 13252 -11338 13286
rect -11372 13184 -11338 13218
rect -11372 13116 -11338 13150
rect -11372 13048 -11338 13082
rect -11372 12980 -11338 13014
rect -11372 12912 -11338 12946
rect -11372 12844 -11338 12878
rect -11372 12776 -11338 12810
rect -11372 12708 -11338 12742
rect -11372 12640 -11338 12674
rect -11372 12572 -11338 12606
rect -11372 12504 -11338 12538
rect -11372 12436 -11338 12470
rect -11372 12368 -11338 12402
rect -11372 12300 -11338 12334
rect -11372 12151 -11338 12266
rect -9016 16516 -8982 16622
rect -9016 16448 -8982 16482
rect -9016 16380 -8982 16414
rect -9016 16312 -8982 16346
rect -9016 16244 -8982 16278
rect -9016 16176 -8982 16210
rect -9016 16108 -8982 16142
rect -9016 16040 -8982 16074
rect -9016 15972 -8982 16006
rect -9016 15904 -8982 15938
rect -9016 15836 -8982 15870
rect -9016 15768 -8982 15802
rect -9016 15700 -8982 15734
rect -9016 15632 -8982 15666
rect -9016 15564 -8982 15598
rect -9016 15496 -8982 15530
rect -9016 15428 -8982 15462
rect -9016 15360 -8982 15394
rect -9016 15292 -8982 15326
rect -9016 15224 -8982 15258
rect -9016 15156 -8982 15190
rect -9016 15088 -8982 15122
rect -9016 15020 -8982 15054
rect -9016 14952 -8982 14986
rect -9016 14884 -8982 14918
rect -9016 14816 -8982 14850
rect -9016 14748 -8982 14782
rect -9016 14680 -8982 14714
rect -9016 14612 -8982 14646
rect -9016 14544 -8982 14578
rect -9016 14476 -8982 14510
rect -9016 14408 -8982 14442
rect -9016 14340 -8982 14374
rect -9016 14272 -8982 14306
rect -9016 14204 -8982 14238
rect -9016 14136 -8982 14170
rect -9016 14068 -8982 14102
rect -9016 14000 -8982 14034
rect -9016 13932 -8982 13966
rect -9016 13864 -8982 13898
rect -9016 13796 -8982 13830
rect -9016 13728 -8982 13762
rect -9016 13660 -8982 13694
rect -9016 13592 -8982 13626
rect -9016 13524 -8982 13558
rect -9016 13456 -8982 13490
rect -9016 13388 -8982 13422
rect -9016 13320 -8982 13354
rect -9016 13252 -8982 13286
rect -9016 13184 -8982 13218
rect -9016 13116 -8982 13150
rect -9016 13048 -8982 13082
rect -9016 12980 -8982 13014
rect -9016 12912 -8982 12946
rect -9016 12844 -8982 12878
rect -9016 12776 -8982 12810
rect -9016 12708 -8982 12742
rect -9016 12640 -8982 12674
rect -9016 12572 -8982 12606
rect -9016 12504 -8982 12538
rect -9016 12436 -8982 12470
rect -9016 12368 -8982 12402
rect -9016 12300 -8982 12334
rect -9016 12151 -8982 12266
rect -11372 12117 -11232 12151
rect -11198 12117 -11164 12151
rect -11130 12117 -11096 12151
rect -11062 12117 -11028 12151
rect -10994 12117 -10960 12151
rect -10926 12117 -10892 12151
rect -10858 12117 -10824 12151
rect -10790 12117 -10756 12151
rect -10722 12117 -10688 12151
rect -10654 12117 -10620 12151
rect -10586 12117 -10552 12151
rect -10518 12117 -10484 12151
rect -10450 12117 -10416 12151
rect -10382 12117 -10348 12151
rect -10314 12117 -10280 12151
rect -10246 12117 -10212 12151
rect -10178 12117 -10144 12151
rect -10110 12117 -10076 12151
rect -10042 12117 -10008 12151
rect -9974 12117 -9940 12151
rect -9906 12117 -9872 12151
rect -9838 12117 -9804 12151
rect -9770 12117 -9736 12151
rect -9702 12117 -9668 12151
rect -9634 12117 -9600 12151
rect -9566 12117 -9532 12151
rect -9498 12117 -9464 12151
rect -9430 12117 -9396 12151
rect -9362 12117 -9328 12151
rect -9294 12117 -9260 12151
rect -9226 12117 -9192 12151
rect -9158 12117 -8982 12151
<< nsubdiffcont >>
rect -11285 16622 -11251 16656
rect -11217 16622 -11183 16656
rect -11149 16622 -11115 16656
rect -11081 16622 -11047 16656
rect -11013 16622 -10979 16656
rect -10945 16622 -10911 16656
rect -10877 16622 -10843 16656
rect -10809 16622 -10775 16656
rect -10741 16622 -10707 16656
rect -10673 16622 -10639 16656
rect -10605 16622 -10571 16656
rect -10537 16622 -10503 16656
rect -10469 16622 -10435 16656
rect -10401 16622 -10367 16656
rect -10333 16622 -10299 16656
rect -10265 16622 -10231 16656
rect -10197 16622 -10163 16656
rect -10129 16622 -10095 16656
rect -10061 16622 -10027 16656
rect -9993 16622 -9959 16656
rect -9925 16622 -9891 16656
rect -9857 16622 -9823 16656
rect -9789 16622 -9755 16656
rect -9721 16622 -9687 16656
rect -9653 16622 -9619 16656
rect -9585 16622 -9551 16656
rect -9517 16622 -9483 16656
rect -9449 16622 -9415 16656
rect -9381 16622 -9347 16656
rect -9313 16622 -9279 16656
rect -9245 16622 -9211 16656
rect -9177 16622 -9143 16656
rect -11372 16482 -11338 16516
rect -11372 16414 -11338 16448
rect -11372 16346 -11338 16380
rect -11372 16278 -11338 16312
rect -11372 16210 -11338 16244
rect -11372 16142 -11338 16176
rect -11372 16074 -11338 16108
rect -11372 16006 -11338 16040
rect -11372 15938 -11338 15972
rect -11372 15870 -11338 15904
rect -11372 15802 -11338 15836
rect -11372 15734 -11338 15768
rect -11372 15666 -11338 15700
rect -11372 15598 -11338 15632
rect -11372 15530 -11338 15564
rect -11372 15462 -11338 15496
rect -11372 15394 -11338 15428
rect -11372 15326 -11338 15360
rect -11372 15258 -11338 15292
rect -11372 15190 -11338 15224
rect -11372 15122 -11338 15156
rect -11372 15054 -11338 15088
rect -11372 14986 -11338 15020
rect -11372 14918 -11338 14952
rect -11372 14850 -11338 14884
rect -11372 14782 -11338 14816
rect -11372 14714 -11338 14748
rect -11372 14646 -11338 14680
rect -11372 14578 -11338 14612
rect -11372 14510 -11338 14544
rect -11372 14442 -11338 14476
rect -11372 14374 -11338 14408
rect -11372 14306 -11338 14340
rect -11372 14238 -11338 14272
rect -11372 14170 -11338 14204
rect -11372 14102 -11338 14136
rect -11372 14034 -11338 14068
rect -11372 13966 -11338 14000
rect -11372 13898 -11338 13932
rect -11372 13830 -11338 13864
rect -11372 13762 -11338 13796
rect -11372 13694 -11338 13728
rect -11372 13626 -11338 13660
rect -11372 13558 -11338 13592
rect -11372 13490 -11338 13524
rect -11372 13422 -11338 13456
rect -11372 13354 -11338 13388
rect -11372 13286 -11338 13320
rect -11372 13218 -11338 13252
rect -11372 13150 -11338 13184
rect -11372 13082 -11338 13116
rect -11372 13014 -11338 13048
rect -11372 12946 -11338 12980
rect -11372 12878 -11338 12912
rect -11372 12810 -11338 12844
rect -11372 12742 -11338 12776
rect -11372 12674 -11338 12708
rect -11372 12606 -11338 12640
rect -11372 12538 -11338 12572
rect -11372 12470 -11338 12504
rect -11372 12402 -11338 12436
rect -11372 12334 -11338 12368
rect -11372 12266 -11338 12300
rect -9016 16482 -8982 16516
rect -9016 16414 -8982 16448
rect -9016 16346 -8982 16380
rect -9016 16278 -8982 16312
rect -9016 16210 -8982 16244
rect -9016 16142 -8982 16176
rect -9016 16074 -8982 16108
rect -9016 16006 -8982 16040
rect -9016 15938 -8982 15972
rect -9016 15870 -8982 15904
rect -9016 15802 -8982 15836
rect -9016 15734 -8982 15768
rect -9016 15666 -8982 15700
rect -9016 15598 -8982 15632
rect -9016 15530 -8982 15564
rect -9016 15462 -8982 15496
rect -9016 15394 -8982 15428
rect -9016 15326 -8982 15360
rect -9016 15258 -8982 15292
rect -9016 15190 -8982 15224
rect -9016 15122 -8982 15156
rect -9016 15054 -8982 15088
rect -9016 14986 -8982 15020
rect -9016 14918 -8982 14952
rect -9016 14850 -8982 14884
rect -9016 14782 -8982 14816
rect -9016 14714 -8982 14748
rect -9016 14646 -8982 14680
rect -9016 14578 -8982 14612
rect -9016 14510 -8982 14544
rect -9016 14442 -8982 14476
rect -9016 14374 -8982 14408
rect -9016 14306 -8982 14340
rect -9016 14238 -8982 14272
rect -9016 14170 -8982 14204
rect -9016 14102 -8982 14136
rect -9016 14034 -8982 14068
rect -9016 13966 -8982 14000
rect -9016 13898 -8982 13932
rect -9016 13830 -8982 13864
rect -9016 13762 -8982 13796
rect -9016 13694 -8982 13728
rect -9016 13626 -8982 13660
rect -9016 13558 -8982 13592
rect -9016 13490 -8982 13524
rect -9016 13422 -8982 13456
rect -9016 13354 -8982 13388
rect -9016 13286 -8982 13320
rect -9016 13218 -8982 13252
rect -9016 13150 -8982 13184
rect -9016 13082 -8982 13116
rect -9016 13014 -8982 13048
rect -9016 12946 -8982 12980
rect -9016 12878 -8982 12912
rect -9016 12810 -8982 12844
rect -9016 12742 -8982 12776
rect -9016 12674 -8982 12708
rect -9016 12606 -8982 12640
rect -9016 12538 -8982 12572
rect -9016 12470 -8982 12504
rect -9016 12402 -8982 12436
rect -9016 12334 -8982 12368
rect -9016 12266 -8982 12300
rect -11232 12117 -11198 12151
rect -11164 12117 -11130 12151
rect -11096 12117 -11062 12151
rect -11028 12117 -10994 12151
rect -10960 12117 -10926 12151
rect -10892 12117 -10858 12151
rect -10824 12117 -10790 12151
rect -10756 12117 -10722 12151
rect -10688 12117 -10654 12151
rect -10620 12117 -10586 12151
rect -10552 12117 -10518 12151
rect -10484 12117 -10450 12151
rect -10416 12117 -10382 12151
rect -10348 12117 -10314 12151
rect -10280 12117 -10246 12151
rect -10212 12117 -10178 12151
rect -10144 12117 -10110 12151
rect -10076 12117 -10042 12151
rect -10008 12117 -9974 12151
rect -9940 12117 -9906 12151
rect -9872 12117 -9838 12151
rect -9804 12117 -9770 12151
rect -9736 12117 -9702 12151
rect -9668 12117 -9634 12151
rect -9600 12117 -9566 12151
rect -9532 12117 -9498 12151
rect -9464 12117 -9430 12151
rect -9396 12117 -9362 12151
rect -9328 12117 -9294 12151
rect -9260 12117 -9226 12151
rect -9192 12117 -9158 12151
<< locali >>
rect -11372 16622 -11285 16656
rect -11251 16622 -11217 16656
rect -11183 16622 -11149 16656
rect -11115 16622 -11081 16656
rect -11047 16622 -11013 16656
rect -10979 16622 -10945 16656
rect -10911 16622 -10877 16656
rect -10843 16622 -10809 16656
rect -10775 16622 -10741 16656
rect -10707 16622 -10673 16656
rect -10639 16622 -10605 16656
rect -10571 16622 -10537 16656
rect -10503 16622 -10469 16656
rect -10435 16622 -10401 16656
rect -10367 16622 -10333 16656
rect -10299 16622 -10265 16656
rect -10231 16622 -10197 16656
rect -10163 16622 -10129 16656
rect -10095 16622 -10061 16656
rect -10027 16622 -9993 16656
rect -9959 16622 -9925 16656
rect -9891 16622 -9857 16656
rect -9823 16622 -9789 16656
rect -9755 16622 -9721 16656
rect -9687 16622 -9653 16656
rect -9619 16622 -9585 16656
rect -9551 16622 -9517 16656
rect -9483 16622 -9449 16656
rect -9415 16622 -9381 16656
rect -9347 16622 -9313 16656
rect -9279 16622 -9245 16656
rect -9211 16622 -9177 16656
rect -9143 16622 -8982 16656
rect -11372 16516 -11338 16622
rect -11372 16448 -11338 16482
rect -11372 16380 -11338 16414
rect -11372 16312 -11338 16346
rect -11372 16244 -11338 16278
rect -11372 16176 -11338 16210
rect -11372 16108 -11338 16142
rect -11372 16040 -11338 16074
rect -11372 15972 -11338 16006
rect -11372 15904 -11338 15938
rect -11372 15836 -11338 15870
rect -11372 15768 -11338 15802
rect -11372 15700 -11338 15734
rect -11372 15632 -11338 15666
rect -11372 15564 -11338 15598
rect -11372 15496 -11338 15530
rect -11372 15428 -11338 15462
rect -11372 15360 -11338 15394
rect -11372 15292 -11338 15326
rect -11372 15224 -11338 15258
rect -11372 15156 -11338 15190
rect -11372 15088 -11338 15122
rect -11372 15020 -11338 15054
rect -11372 14952 -11338 14986
rect -11372 14884 -11338 14918
rect -11372 14816 -11338 14850
rect -11372 14748 -11338 14782
rect -11372 14680 -11338 14714
rect -11372 14612 -11338 14646
rect -11372 14544 -11338 14578
rect -11372 14476 -11338 14510
rect -11372 14408 -11338 14442
rect -11372 14340 -11338 14374
rect -11372 14272 -11338 14306
rect -11372 14204 -11338 14238
rect -11372 14136 -11338 14170
rect -11372 14068 -11338 14102
rect -11372 14000 -11338 14034
rect -11372 13932 -11338 13966
rect -11372 13864 -11338 13898
rect -11372 13796 -11338 13830
rect -11372 13728 -11338 13762
rect -11372 13660 -11338 13694
rect -11372 13592 -11338 13626
rect -11372 13524 -11338 13558
rect -11372 13456 -11338 13490
rect -11372 13388 -11338 13422
rect -11372 13320 -11338 13354
rect -11372 13252 -11338 13286
rect -11372 13184 -11338 13218
rect -11372 13116 -11338 13150
rect -11372 13048 -11338 13082
rect -11372 12980 -11338 13014
rect -11372 12912 -11338 12946
rect -11372 12844 -11338 12878
rect -11372 12776 -11338 12810
rect -11372 12708 -11338 12742
rect -11372 12640 -11338 12674
rect -11372 12572 -11338 12606
rect -11372 12504 -11338 12538
rect -11372 12436 -11338 12470
rect -11372 12368 -11338 12402
rect -11372 12300 -11338 12334
rect -11372 12151 -11338 12266
rect -9016 16516 -8982 16622
rect -9016 16448 -8982 16482
rect -9016 16380 -8982 16414
rect -9016 16312 -8982 16346
rect -9016 16244 -8982 16278
rect -9016 16176 -8982 16210
rect -9016 16108 -8982 16142
rect -9016 16040 -8982 16074
rect -9016 15972 -8982 16006
rect -9016 15904 -8982 15938
rect -9016 15836 -8982 15870
rect -9016 15768 -8982 15802
rect -9016 15700 -8982 15734
rect -9016 15632 -8982 15666
rect -9016 15564 -8982 15598
rect -9016 15496 -8982 15530
rect -9016 15428 -8982 15462
rect -9016 15360 -8982 15394
rect -9016 15292 -8982 15326
rect -9016 15224 -8982 15258
rect -9016 15156 -8982 15190
rect -9016 15088 -8982 15122
rect -9016 15020 -8982 15054
rect -9016 14952 -8982 14986
rect -9016 14884 -8982 14918
rect -9016 14816 -8982 14850
rect -9016 14748 -8982 14782
rect -9016 14680 -8982 14714
rect -9016 14612 -8982 14646
rect -9016 14544 -8982 14578
rect -9016 14476 -8982 14510
rect -9016 14408 -8982 14442
rect -9016 14340 -8982 14374
rect -9016 14272 -8982 14306
rect -9016 14204 -8982 14238
rect -9016 14136 -8982 14170
rect -9016 14068 -8982 14102
rect -9016 14000 -8982 14034
rect -9016 13932 -8982 13966
rect -9016 13864 -8982 13898
rect -9016 13796 -8982 13830
rect -9016 13728 -8982 13762
rect -9016 13660 -8982 13694
rect -9016 13592 -8982 13626
rect -9016 13524 -8982 13558
rect -9016 13456 -8982 13490
rect -9016 13388 -8982 13422
rect -9016 13320 -8982 13354
rect -9016 13252 -8982 13286
rect -9016 13184 -8982 13218
rect -9016 13116 -8982 13150
rect -9016 13048 -8982 13082
rect -9016 12980 -8982 13014
rect -9016 12912 -8982 12946
rect -9016 12844 -8982 12878
rect -9016 12776 -8982 12810
rect -9016 12708 -8982 12742
rect -9016 12640 -8982 12674
rect -9016 12572 -8982 12606
rect -9016 12504 -8982 12538
rect -9016 12436 -8982 12470
rect -9016 12368 -8982 12402
rect -9016 12300 -8982 12334
rect -9016 12151 -8982 12266
rect -11372 12117 -11232 12151
rect -11198 12117 -11164 12151
rect -11130 12117 -11096 12151
rect -11062 12117 -11028 12151
rect -10994 12117 -10960 12151
rect -10926 12117 -10892 12151
rect -10858 12117 -10824 12151
rect -10790 12117 -10756 12151
rect -10722 12117 -10688 12151
rect -10654 12117 -10620 12151
rect -10586 12117 -10552 12151
rect -10518 12117 -10484 12151
rect -10450 12117 -10416 12151
rect -10382 12117 -10348 12151
rect -10314 12117 -10280 12151
rect -10246 12117 -10212 12151
rect -10178 12117 -10144 12151
rect -10110 12117 -10076 12151
rect -10042 12117 -10008 12151
rect -9974 12117 -9940 12151
rect -9906 12117 -9872 12151
rect -9838 12117 -9804 12151
rect -9770 12117 -9736 12151
rect -9702 12117 -9668 12151
rect -9634 12117 -9600 12151
rect -9566 12117 -9532 12151
rect -9498 12117 -9464 12151
rect -9430 12117 -9396 12151
rect -9362 12117 -9328 12151
rect -9294 12117 -9260 12151
rect -9226 12117 -9192 12151
rect -9158 12117 -8982 12151
<< properties >>
string path -57.040 83.195 -44.995 83.195 -44.995 60.670 -56.775 60.670 -56.775 83.195 
<< end >>
