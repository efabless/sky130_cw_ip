magic
tech sky130A
magscale 1 2
timestamp 1715010268
<< pwell >>
rect -350 1202 350 1288
rect -350 -1202 -264 1202
rect 264 -1202 350 1202
rect -350 -1288 350 -1202
<< psubdiff >>
rect -324 1228 -221 1262
rect -187 1228 -153 1262
rect -119 1228 -85 1262
rect -51 1228 -17 1262
rect 17 1228 51 1262
rect 85 1228 119 1262
rect 153 1228 187 1262
rect 221 1228 324 1262
rect -324 1139 -290 1228
rect 290 1139 324 1228
rect -324 1071 -290 1105
rect -324 1003 -290 1037
rect -324 935 -290 969
rect -324 867 -290 901
rect -324 799 -290 833
rect -324 731 -290 765
rect -324 663 -290 697
rect -324 595 -290 629
rect -324 527 -290 561
rect -324 459 -290 493
rect -324 391 -290 425
rect -324 323 -290 357
rect -324 255 -290 289
rect -324 187 -290 221
rect -324 119 -290 153
rect -324 51 -290 85
rect -324 -17 -290 17
rect -324 -85 -290 -51
rect -324 -153 -290 -119
rect -324 -221 -290 -187
rect -324 -289 -290 -255
rect -324 -357 -290 -323
rect -324 -425 -290 -391
rect -324 -493 -290 -459
rect -324 -561 -290 -527
rect -324 -629 -290 -595
rect -324 -697 -290 -663
rect -324 -765 -290 -731
rect -324 -833 -290 -799
rect -324 -901 -290 -867
rect -324 -969 -290 -935
rect -324 -1037 -290 -1003
rect -324 -1105 -290 -1071
rect 290 1071 324 1105
rect 290 1003 324 1037
rect 290 935 324 969
rect 290 867 324 901
rect 290 799 324 833
rect 290 731 324 765
rect 290 663 324 697
rect 290 595 324 629
rect 290 527 324 561
rect 290 459 324 493
rect 290 391 324 425
rect 290 323 324 357
rect 290 255 324 289
rect 290 187 324 221
rect 290 119 324 153
rect 290 51 324 85
rect 290 -17 324 17
rect 290 -85 324 -51
rect 290 -153 324 -119
rect 290 -221 324 -187
rect 290 -289 324 -255
rect 290 -357 324 -323
rect 290 -425 324 -391
rect 290 -493 324 -459
rect 290 -561 324 -527
rect 290 -629 324 -595
rect 290 -697 324 -663
rect 290 -765 324 -731
rect 290 -833 324 -799
rect 290 -901 324 -867
rect 290 -969 324 -935
rect 290 -1037 324 -1003
rect 290 -1105 324 -1071
rect -324 -1228 -290 -1139
rect 290 -1228 324 -1139
rect -324 -1262 -221 -1228
rect -187 -1262 -153 -1228
rect -119 -1262 -85 -1228
rect -51 -1262 -17 -1228
rect 17 -1262 51 -1228
rect 85 -1262 119 -1228
rect 153 -1262 187 -1228
rect 221 -1262 324 -1228
<< psubdiffcont >>
rect -221 1228 -187 1262
rect -153 1228 -119 1262
rect -85 1228 -51 1262
rect -17 1228 17 1262
rect 51 1228 85 1262
rect 119 1228 153 1262
rect 187 1228 221 1262
rect -324 1105 -290 1139
rect -324 1037 -290 1071
rect -324 969 -290 1003
rect -324 901 -290 935
rect -324 833 -290 867
rect -324 765 -290 799
rect -324 697 -290 731
rect -324 629 -290 663
rect -324 561 -290 595
rect -324 493 -290 527
rect -324 425 -290 459
rect -324 357 -290 391
rect -324 289 -290 323
rect -324 221 -290 255
rect -324 153 -290 187
rect -324 85 -290 119
rect -324 17 -290 51
rect -324 -51 -290 -17
rect -324 -119 -290 -85
rect -324 -187 -290 -153
rect -324 -255 -290 -221
rect -324 -323 -290 -289
rect -324 -391 -290 -357
rect -324 -459 -290 -425
rect -324 -527 -290 -493
rect -324 -595 -290 -561
rect -324 -663 -290 -629
rect -324 -731 -290 -697
rect -324 -799 -290 -765
rect -324 -867 -290 -833
rect -324 -935 -290 -901
rect -324 -1003 -290 -969
rect -324 -1071 -290 -1037
rect -324 -1139 -290 -1105
rect 290 1105 324 1139
rect 290 1037 324 1071
rect 290 969 324 1003
rect 290 901 324 935
rect 290 833 324 867
rect 290 765 324 799
rect 290 697 324 731
rect 290 629 324 663
rect 290 561 324 595
rect 290 493 324 527
rect 290 425 324 459
rect 290 357 324 391
rect 290 289 324 323
rect 290 221 324 255
rect 290 153 324 187
rect 290 85 324 119
rect 290 17 324 51
rect 290 -51 324 -17
rect 290 -119 324 -85
rect 290 -187 324 -153
rect 290 -255 324 -221
rect 290 -323 324 -289
rect 290 -391 324 -357
rect 290 -459 324 -425
rect 290 -527 324 -493
rect 290 -595 324 -561
rect 290 -663 324 -629
rect 290 -731 324 -697
rect 290 -799 324 -765
rect 290 -867 324 -833
rect 290 -935 324 -901
rect 290 -1003 324 -969
rect 290 -1071 324 -1037
rect 290 -1139 324 -1105
rect -221 -1262 -187 -1228
rect -153 -1262 -119 -1228
rect -85 -1262 -51 -1228
rect -17 -1262 17 -1228
rect 51 -1262 85 -1228
rect 119 -1262 153 -1228
rect 187 -1262 221 -1228
<< xpolycontact >>
rect -194 696 -124 1132
rect -194 -1132 -124 -696
rect 124 696 194 1132
rect 124 -1132 194 -696
<< xpolyres >>
rect -194 -696 -124 696
rect 124 -696 194 696
<< locali >>
rect -324 1228 -221 1262
rect -187 1228 -153 1262
rect -119 1228 -85 1262
rect -51 1228 -17 1262
rect 17 1228 51 1262
rect 85 1228 119 1262
rect 153 1228 187 1262
rect 221 1228 324 1262
rect -324 1139 -290 1228
rect 290 1139 324 1228
rect -324 1071 -290 1105
rect -324 1003 -290 1037
rect -324 935 -290 969
rect -324 867 -290 901
rect -324 799 -290 833
rect -324 731 -290 765
rect -324 663 -290 697
rect 290 1071 324 1105
rect 290 1003 324 1037
rect 290 935 324 969
rect 290 867 324 901
rect 290 799 324 833
rect 290 731 324 765
rect -324 595 -290 629
rect -324 527 -290 561
rect -324 459 -290 493
rect -324 391 -290 425
rect -324 323 -290 357
rect -324 255 -290 289
rect -324 187 -290 221
rect -324 119 -290 153
rect -324 51 -290 85
rect -324 -17 -290 17
rect -324 -85 -290 -51
rect -324 -153 -290 -119
rect -324 -221 -290 -187
rect -324 -289 -290 -255
rect -324 -357 -290 -323
rect -324 -425 -290 -391
rect -324 -493 -290 -459
rect -324 -561 -290 -527
rect -324 -629 -290 -595
rect -324 -697 -290 -663
rect 290 663 324 697
rect 290 595 324 629
rect 290 527 324 561
rect 290 459 324 493
rect 290 391 324 425
rect 290 323 324 357
rect 290 255 324 289
rect 290 187 324 221
rect 290 119 324 153
rect 290 51 324 85
rect 290 -17 324 17
rect 290 -85 324 -51
rect 290 -153 324 -119
rect 290 -221 324 -187
rect 290 -289 324 -255
rect 290 -357 324 -323
rect 290 -425 324 -391
rect 290 -493 324 -459
rect 290 -561 324 -527
rect 290 -629 324 -595
rect -324 -765 -290 -731
rect -324 -833 -290 -799
rect -324 -901 -290 -867
rect -324 -969 -290 -935
rect -324 -1037 -290 -1003
rect -324 -1105 -290 -1071
rect 290 -697 324 -663
rect 290 -765 324 -731
rect 290 -833 324 -799
rect 290 -901 324 -867
rect 290 -969 324 -935
rect 290 -1037 324 -1003
rect 290 -1105 324 -1071
rect -324 -1228 -290 -1139
rect 290 -1228 324 -1139
rect -324 -1262 -221 -1228
rect -187 -1262 -153 -1228
rect -119 -1262 -85 -1228
rect -51 -1262 -17 -1228
rect 17 -1262 51 -1228
rect 85 -1262 119 -1228
rect 153 -1262 187 -1228
rect 221 -1262 324 -1228
<< viali >>
rect -176 1078 -142 1112
rect -176 1006 -142 1040
rect -176 934 -142 968
rect -176 862 -142 896
rect -176 790 -142 824
rect -176 718 -142 752
rect 142 1078 176 1112
rect 142 1006 176 1040
rect 142 934 176 968
rect 142 862 176 896
rect 142 790 176 824
rect 142 718 176 752
rect -176 -753 -142 -719
rect -176 -825 -142 -791
rect -176 -897 -142 -863
rect -176 -969 -142 -935
rect -176 -1041 -142 -1007
rect -176 -1113 -142 -1079
rect 142 -753 176 -719
rect 142 -825 176 -791
rect 142 -897 176 -863
rect 142 -969 176 -935
rect 142 -1041 176 -1007
rect 142 -1113 176 -1079
<< metal1 >>
rect -184 1112 -134 1126
rect -184 1078 -176 1112
rect -142 1078 -134 1112
rect -184 1040 -134 1078
rect -184 1006 -176 1040
rect -142 1006 -134 1040
rect -184 968 -134 1006
rect -184 934 -176 968
rect -142 934 -134 968
rect -184 896 -134 934
rect -184 862 -176 896
rect -142 862 -134 896
rect -184 824 -134 862
rect -184 790 -176 824
rect -142 790 -134 824
rect -184 752 -134 790
rect -184 718 -176 752
rect -142 718 -134 752
rect -184 705 -134 718
rect 134 1112 184 1126
rect 134 1078 142 1112
rect 176 1078 184 1112
rect 134 1040 184 1078
rect 134 1006 142 1040
rect 176 1006 184 1040
rect 134 968 184 1006
rect 134 934 142 968
rect 176 934 184 968
rect 134 896 184 934
rect 134 862 142 896
rect 176 862 184 896
rect 134 824 184 862
rect 134 790 142 824
rect 176 790 184 824
rect 134 752 184 790
rect 134 718 142 752
rect 176 718 184 752
rect 134 705 184 718
rect -184 -719 -134 -705
rect -184 -753 -176 -719
rect -142 -753 -134 -719
rect -184 -791 -134 -753
rect -184 -825 -176 -791
rect -142 -825 -134 -791
rect -184 -863 -134 -825
rect -184 -897 -176 -863
rect -142 -897 -134 -863
rect -184 -935 -134 -897
rect -184 -969 -176 -935
rect -142 -969 -134 -935
rect -184 -1007 -134 -969
rect -184 -1041 -176 -1007
rect -142 -1041 -134 -1007
rect -184 -1079 -134 -1041
rect -184 -1113 -176 -1079
rect -142 -1113 -134 -1079
rect -184 -1126 -134 -1113
rect 134 -719 184 -705
rect 134 -753 142 -719
rect 176 -753 184 -719
rect 134 -791 184 -753
rect 134 -825 142 -791
rect 176 -825 184 -791
rect 134 -863 184 -825
rect 134 -897 142 -863
rect 176 -897 184 -863
rect 134 -935 184 -897
rect 134 -969 142 -935
rect 176 -969 184 -935
rect 134 -1007 184 -969
rect 134 -1041 142 -1007
rect 176 -1041 184 -1007
rect 134 -1079 184 -1041
rect 134 -1113 142 -1079
rect 176 -1113 184 -1079
rect 134 -1126 184 -1113
<< properties >>
string FIXED_BBOX -307 -1245 307 1245
<< end >>
