magic
tech sky130A
magscale 1 2
timestamp 1715010268
<< pwell >>
rect -273 2419 2505 2505
rect -273 -187 -187 2419
rect 2419 -187 2505 2419
rect -273 -273 2505 -187
<< psubdiff >>
rect -247 2445 -67 2479
rect -33 2445 1 2479
rect 35 2445 69 2479
rect 103 2445 137 2479
rect 171 2445 205 2479
rect 239 2445 273 2479
rect 307 2445 341 2479
rect 375 2445 409 2479
rect 443 2445 477 2479
rect 511 2445 545 2479
rect 579 2445 613 2479
rect 647 2445 681 2479
rect 715 2445 749 2479
rect 783 2445 817 2479
rect 851 2445 885 2479
rect 919 2445 953 2479
rect 987 2445 1021 2479
rect 1055 2445 1089 2479
rect 1123 2445 1157 2479
rect 1191 2445 1225 2479
rect 1259 2445 1293 2479
rect 1327 2445 1361 2479
rect 1395 2445 1429 2479
rect 1463 2445 1497 2479
rect 1531 2445 1565 2479
rect 1599 2445 1633 2479
rect 1667 2445 1701 2479
rect 1735 2445 1769 2479
rect 1803 2445 1837 2479
rect 1871 2445 1905 2479
rect 1939 2445 1973 2479
rect 2007 2445 2041 2479
rect 2075 2445 2109 2479
rect 2143 2445 2177 2479
rect 2211 2445 2245 2479
rect 2279 2445 2479 2479
rect -247 2279 -213 2445
rect -247 2211 -213 2245
rect -247 2143 -213 2177
rect -247 2075 -213 2109
rect -247 2007 -213 2041
rect -247 1939 -213 1973
rect -247 1871 -213 1905
rect -247 1803 -213 1837
rect -247 1735 -213 1769
rect -247 1667 -213 1701
rect -247 1599 -213 1633
rect -247 1531 -213 1565
rect -247 1463 -213 1497
rect -247 1395 -213 1429
rect -247 1327 -213 1361
rect -247 1259 -213 1293
rect -247 1191 -213 1225
rect -247 1123 -213 1157
rect -247 1055 -213 1089
rect -247 987 -213 1021
rect -247 919 -213 953
rect -247 851 -213 885
rect -247 783 -213 817
rect -247 715 -213 749
rect -247 647 -213 681
rect -247 579 -213 613
rect -247 511 -213 545
rect -247 443 -213 477
rect -247 375 -213 409
rect -247 307 -213 341
rect -247 239 -213 273
rect -247 171 -213 205
rect -247 103 -213 137
rect -247 35 -213 69
rect -247 -213 -213 1
rect 2445 2279 2479 2445
rect 2445 2211 2479 2245
rect 2445 2143 2479 2177
rect 2445 2075 2479 2109
rect 2445 2007 2479 2041
rect 2445 1939 2479 1973
rect 2445 1871 2479 1905
rect 2445 1803 2479 1837
rect 2445 1735 2479 1769
rect 2445 1667 2479 1701
rect 2445 1599 2479 1633
rect 2445 1531 2479 1565
rect 2445 1463 2479 1497
rect 2445 1395 2479 1429
rect 2445 1327 2479 1361
rect 2445 1259 2479 1293
rect 2445 1191 2479 1225
rect 2445 1123 2479 1157
rect 2445 1055 2479 1089
rect 2445 987 2479 1021
rect 2445 919 2479 953
rect 2445 851 2479 885
rect 2445 783 2479 817
rect 2445 715 2479 749
rect 2445 647 2479 681
rect 2445 579 2479 613
rect 2445 511 2479 545
rect 2445 443 2479 477
rect 2445 375 2479 409
rect 2445 307 2479 341
rect 2445 239 2479 273
rect 2445 171 2479 205
rect 2445 103 2479 137
rect 2445 35 2479 69
rect 2445 -213 2479 1
rect -247 -247 1 -213
rect 35 -247 69 -213
rect 103 -247 137 -213
rect 171 -247 205 -213
rect 239 -247 273 -213
rect 307 -247 341 -213
rect 375 -247 409 -213
rect 443 -247 477 -213
rect 511 -247 545 -213
rect 579 -247 613 -213
rect 647 -247 681 -213
rect 715 -247 749 -213
rect 783 -247 817 -213
rect 851 -247 885 -213
rect 919 -247 953 -213
rect 987 -247 1021 -213
rect 1055 -247 1089 -213
rect 1123 -247 1157 -213
rect 1191 -247 1225 -213
rect 1259 -247 1293 -213
rect 1327 -247 1361 -213
rect 1395 -247 1429 -213
rect 1463 -247 1497 -213
rect 1531 -247 1565 -213
rect 1599 -247 1633 -213
rect 1667 -247 1701 -213
rect 1735 -247 1769 -213
rect 1803 -247 1837 -213
rect 1871 -247 1905 -213
rect 1939 -247 1973 -213
rect 2007 -247 2041 -213
rect 2075 -247 2109 -213
rect 2143 -247 2177 -213
rect 2211 -247 2245 -213
rect 2279 -247 2479 -213
<< psubdiffcont >>
rect -67 2445 -33 2479
rect 1 2445 35 2479
rect 69 2445 103 2479
rect 137 2445 171 2479
rect 205 2445 239 2479
rect 273 2445 307 2479
rect 341 2445 375 2479
rect 409 2445 443 2479
rect 477 2445 511 2479
rect 545 2445 579 2479
rect 613 2445 647 2479
rect 681 2445 715 2479
rect 749 2445 783 2479
rect 817 2445 851 2479
rect 885 2445 919 2479
rect 953 2445 987 2479
rect 1021 2445 1055 2479
rect 1089 2445 1123 2479
rect 1157 2445 1191 2479
rect 1225 2445 1259 2479
rect 1293 2445 1327 2479
rect 1361 2445 1395 2479
rect 1429 2445 1463 2479
rect 1497 2445 1531 2479
rect 1565 2445 1599 2479
rect 1633 2445 1667 2479
rect 1701 2445 1735 2479
rect 1769 2445 1803 2479
rect 1837 2445 1871 2479
rect 1905 2445 1939 2479
rect 1973 2445 2007 2479
rect 2041 2445 2075 2479
rect 2109 2445 2143 2479
rect 2177 2445 2211 2479
rect 2245 2445 2279 2479
rect -247 2245 -213 2279
rect -247 2177 -213 2211
rect -247 2109 -213 2143
rect -247 2041 -213 2075
rect -247 1973 -213 2007
rect -247 1905 -213 1939
rect -247 1837 -213 1871
rect -247 1769 -213 1803
rect -247 1701 -213 1735
rect -247 1633 -213 1667
rect -247 1565 -213 1599
rect -247 1497 -213 1531
rect -247 1429 -213 1463
rect -247 1361 -213 1395
rect -247 1293 -213 1327
rect -247 1225 -213 1259
rect -247 1157 -213 1191
rect -247 1089 -213 1123
rect -247 1021 -213 1055
rect -247 953 -213 987
rect -247 885 -213 919
rect -247 817 -213 851
rect -247 749 -213 783
rect -247 681 -213 715
rect -247 613 -213 647
rect -247 545 -213 579
rect -247 477 -213 511
rect -247 409 -213 443
rect -247 341 -213 375
rect -247 273 -213 307
rect -247 205 -213 239
rect -247 137 -213 171
rect -247 69 -213 103
rect -247 1 -213 35
rect 2445 2245 2479 2279
rect 2445 2177 2479 2211
rect 2445 2109 2479 2143
rect 2445 2041 2479 2075
rect 2445 1973 2479 2007
rect 2445 1905 2479 1939
rect 2445 1837 2479 1871
rect 2445 1769 2479 1803
rect 2445 1701 2479 1735
rect 2445 1633 2479 1667
rect 2445 1565 2479 1599
rect 2445 1497 2479 1531
rect 2445 1429 2479 1463
rect 2445 1361 2479 1395
rect 2445 1293 2479 1327
rect 2445 1225 2479 1259
rect 2445 1157 2479 1191
rect 2445 1089 2479 1123
rect 2445 1021 2479 1055
rect 2445 953 2479 987
rect 2445 885 2479 919
rect 2445 817 2479 851
rect 2445 749 2479 783
rect 2445 681 2479 715
rect 2445 613 2479 647
rect 2445 545 2479 579
rect 2445 477 2479 511
rect 2445 409 2479 443
rect 2445 341 2479 375
rect 2445 273 2479 307
rect 2445 205 2479 239
rect 2445 137 2479 171
rect 2445 69 2479 103
rect 2445 1 2479 35
rect 1 -247 35 -213
rect 69 -247 103 -213
rect 137 -247 171 -213
rect 205 -247 239 -213
rect 273 -247 307 -213
rect 341 -247 375 -213
rect 409 -247 443 -213
rect 477 -247 511 -213
rect 545 -247 579 -213
rect 613 -247 647 -213
rect 681 -247 715 -213
rect 749 -247 783 -213
rect 817 -247 851 -213
rect 885 -247 919 -213
rect 953 -247 987 -213
rect 1021 -247 1055 -213
rect 1089 -247 1123 -213
rect 1157 -247 1191 -213
rect 1225 -247 1259 -213
rect 1293 -247 1327 -213
rect 1361 -247 1395 -213
rect 1429 -247 1463 -213
rect 1497 -247 1531 -213
rect 1565 -247 1599 -213
rect 1633 -247 1667 -213
rect 1701 -247 1735 -213
rect 1769 -247 1803 -213
rect 1837 -247 1871 -213
rect 1905 -247 1939 -213
rect 1973 -247 2007 -213
rect 2041 -247 2075 -213
rect 2109 -247 2143 -213
rect 2177 -247 2211 -213
rect 2245 -247 2279 -213
<< locali >>
rect -247 2445 -67 2479
rect -33 2445 1 2479
rect 35 2445 69 2479
rect 103 2445 137 2479
rect 171 2445 205 2479
rect 239 2445 273 2479
rect 307 2445 341 2479
rect 375 2445 409 2479
rect 443 2445 477 2479
rect 511 2445 545 2479
rect 579 2445 613 2479
rect 647 2445 681 2479
rect 715 2445 749 2479
rect 783 2445 817 2479
rect 851 2445 885 2479
rect 919 2445 953 2479
rect 987 2445 1021 2479
rect 1055 2445 1089 2479
rect 1123 2445 1157 2479
rect 1191 2445 1225 2479
rect 1259 2445 1293 2479
rect 1327 2445 1361 2479
rect 1395 2445 1429 2479
rect 1463 2445 1497 2479
rect 1531 2445 1565 2479
rect 1599 2445 1633 2479
rect 1667 2445 1701 2479
rect 1735 2445 1769 2479
rect 1803 2445 1837 2479
rect 1871 2445 1905 2479
rect 1939 2445 1973 2479
rect 2007 2445 2041 2479
rect 2075 2445 2109 2479
rect 2143 2445 2177 2479
rect 2211 2445 2245 2479
rect 2279 2445 2479 2479
rect -247 2279 -213 2445
rect -247 2211 -213 2245
rect -247 2143 -213 2177
rect -247 2075 -213 2109
rect -247 2007 -213 2041
rect -247 1939 -213 1973
rect -247 1871 -213 1905
rect -247 1803 -213 1837
rect -247 1735 -213 1769
rect -247 1667 -213 1701
rect -247 1599 -213 1633
rect -247 1531 -213 1565
rect -247 1463 -213 1497
rect -247 1395 -213 1429
rect -247 1327 -213 1361
rect -247 1259 -213 1293
rect -247 1191 -213 1225
rect -247 1123 -213 1157
rect -247 1055 -213 1089
rect -247 987 -213 1021
rect -247 919 -213 953
rect -247 851 -213 885
rect -247 783 -213 817
rect -247 715 -213 749
rect -247 647 -213 681
rect -247 579 -213 613
rect -247 511 -213 545
rect -247 443 -213 477
rect -247 375 -213 409
rect -247 307 -213 341
rect -247 239 -213 273
rect -247 171 -213 205
rect -247 103 -213 137
rect -247 35 -213 69
rect -247 -213 -213 1
rect 2445 2279 2479 2445
rect 2445 2211 2479 2245
rect 2445 2143 2479 2177
rect 2445 2075 2479 2109
rect 2445 2007 2479 2041
rect 2445 1939 2479 1973
rect 2445 1871 2479 1905
rect 2445 1803 2479 1837
rect 2445 1735 2479 1769
rect 2445 1667 2479 1701
rect 2445 1599 2479 1633
rect 2445 1531 2479 1565
rect 2445 1463 2479 1497
rect 2445 1395 2479 1429
rect 2445 1327 2479 1361
rect 2445 1259 2479 1293
rect 2445 1191 2479 1225
rect 2445 1123 2479 1157
rect 2445 1055 2479 1089
rect 2445 987 2479 1021
rect 2445 919 2479 953
rect 2445 851 2479 885
rect 2445 783 2479 817
rect 2445 715 2479 749
rect 2445 647 2479 681
rect 2445 579 2479 613
rect 2445 511 2479 545
rect 2445 443 2479 477
rect 2445 375 2479 409
rect 2445 307 2479 341
rect 2445 239 2479 273
rect 2445 171 2479 205
rect 2445 103 2479 137
rect 2445 35 2479 69
rect 2445 -213 2479 1
rect -247 -247 1 -213
rect 35 -247 69 -213
rect 103 -247 137 -213
rect 171 -247 205 -213
rect 239 -247 273 -213
rect 307 -247 341 -213
rect 375 -247 409 -213
rect 443 -247 477 -213
rect 511 -247 545 -213
rect 579 -247 613 -213
rect 647 -247 681 -213
rect 715 -247 749 -213
rect 783 -247 817 -213
rect 851 -247 885 -213
rect 919 -247 953 -213
rect 987 -247 1021 -213
rect 1055 -247 1089 -213
rect 1123 -247 1157 -213
rect 1191 -247 1225 -213
rect 1259 -247 1293 -213
rect 1327 -247 1361 -213
rect 1395 -247 1429 -213
rect 1463 -247 1497 -213
rect 1531 -247 1565 -213
rect 1599 -247 1633 -213
rect 1667 -247 1701 -213
rect 1735 -247 1769 -213
rect 1803 -247 1837 -213
rect 1871 -247 1905 -213
rect 1939 -247 1973 -213
rect 2007 -247 2041 -213
rect 2075 -247 2109 -213
rect 2143 -247 2177 -213
rect 2211 -247 2245 -213
rect 2279 -247 2479 -213
<< properties >>
string path -6.800 61.550 61.550 61.550 61.550 -5.750 -5.750 -5.750 -5.750 61.550 
<< end >>
