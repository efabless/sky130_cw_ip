magic
tech sky130A
magscale 1 2
timestamp 1715010268
<< poly >>
rect 381 393 581 1824
rect 639 393 839 1824
rect 1055 393 1255 1824
rect 1313 393 1513 1824
rect 1729 393 1929 1824
rect 1987 393 2187 1824
<< metal1 >>
rect 76 2020 2476 2066
rect 76 116 122 2020
rect 234 1768 2239 1814
rect 234 378 280 1768
rect 329 1727 375 1768
rect 845 1727 891 1768
rect 1677 1727 1723 1768
rect 2193 1727 2239 1768
rect 587 445 633 1727
rect 1261 445 1307 1727
rect 1935 445 1981 1727
rect 329 378 375 419
rect 845 378 891 419
rect 1677 378 1723 419
rect 2193 378 2239 419
rect 234 332 2239 378
rect 2430 116 2476 2020
rect 76 70 2476 116
<< metal2 >>
rect 986 1283 1066 1517
rect 1502 1283 1582 1517
rect 59 1112 139 1271
rect 312 1203 2389 1283
rect 59 1032 2008 1112
rect 59 871 139 1032
rect 2309 729 2389 1203
rect 986 649 2389 729
rect 164 0 244 602
rect 2309 0 2389 649
<< metal3 >>
rect 0 1032 298 1112
rect 986 863 2549 943
use bbp__Guardring_P  bbp__Guardring_P_0
timestamp 1715010268
transform 1 0 0 0 1 -30
box 46 70 2506 2126
use bbp__M4  bbp__M4_0
timestamp 1715010268
transform 1 0 1413 0 1 1663
box -194 -198 194 164
use bbp__M4  bbp__M4_1
timestamp 1715010268
transform 1 0 1155 0 1 1663
box -194 -198 194 164
use bbp__M4  bbp__M4_2
timestamp 1715010268
transform 1 0 1155 0 -1 483
box -194 -198 194 164
use bbp__M4  bbp__M4_3
timestamp 1715010268
transform 1 0 1413 0 -1 483
box -194 -198 194 164
use bbp__M4_nc  bbp__M4_nc_0
timestamp 1715010268
transform 1 0 739 0 1 1109
box -194 -198 194 126
use bbp__M4_nc  bbp__M4_nc_1
timestamp 1715010268
transform 1 0 2087 0 1 1109
box -194 -198 194 126
use bbp__M4_nc  bbp__M4_nc_2
timestamp 1715010268
transform 1 0 1829 0 1 1109
box -194 -198 194 126
use bbp__M4_nc  bbp__M4_nc_3
timestamp 1715010268
transform 1 0 481 0 1 1109
box -194 -198 194 126
use bbp__M5  bbp__M5_0
timestamp 1715010268
transform 1 0 2087 0 1 1663
box -194 -198 194 164
use bbp__M5  bbp__M5_1
timestamp 1715010268
transform 1 0 1829 0 1 1663
box -194 -198 194 164
use bbp__M5  bbp__M5_2
timestamp 1715010268
transform 1 0 739 0 1 1663
box -194 -198 194 164
use bbp__M5  bbp__M5_3
timestamp 1715010268
transform 1 0 481 0 -1 483
box -194 -198 194 164
use bbp__M5  bbp__M5_4
timestamp 1715010268
transform 1 0 739 0 -1 483
box -194 -198 194 164
use bbp__M5  bbp__M5_5
timestamp 1715010268
transform 1 0 1829 0 -1 483
box -194 -198 194 164
use bbp__M5  bbp__M5_6
timestamp 1715010268
transform 1 0 2087 0 -1 483
box -194 -198 194 164
use bbp__M5  bbp__M5_7
timestamp 1715010268
transform 1 0 481 0 1 1663
box -194 -198 194 164
use bbp__M6  bbp__M6_0
timestamp 1715010268
transform 1 0 1413 0 1 1109
box -194 -198 194 126
use bbp__M6  bbp__M6_1
timestamp 1715010268
transform 1 0 1155 0 1 1109
box -194 -198 194 126
use via__LI_M1  via__LI_M1_0
timestamp 1715010268
transform 0 -1 2476 1 0 1190
box -6 -6 124 52
use via__LI_M1  via__LI_M1_1
timestamp 1715010268
transform 0 -1 2476 1 0 1390
box -6 -6 124 52
use via__LI_M1  via__LI_M1_2
timestamp 1715010268
transform 0 -1 2476 1 0 1590
box -6 -6 124 52
use via__LI_M1  via__LI_M1_3
timestamp 1715010268
transform 0 -1 2476 1 0 1790
box -6 -6 124 52
use via__LI_M1  via__LI_M1_4
timestamp 1715010268
transform -1 0 2207 0 -1 2066
box -6 -6 124 52
use via__LI_M1  via__LI_M1_5
timestamp 1715010268
transform -1 0 2007 0 -1 2066
box -6 -6 124 52
use via__LI_M1  via__LI_M1_6
timestamp 1715010268
transform -1 0 1807 0 -1 2066
box -6 -6 124 52
use via__LI_M1  via__LI_M1_7
timestamp 1715010268
transform -1 0 1607 0 -1 2066
box -6 -6 124 52
use via__LI_M1  via__LI_M1_8
timestamp 1715010268
transform -1 0 1407 0 -1 2066
box -6 -6 124 52
use via__LI_M1  via__LI_M1_9
timestamp 1715010268
transform -1 0 1207 0 -1 2066
box -6 -6 124 52
use via__LI_M1  via__LI_M1_10
timestamp 1715010268
transform -1 0 1007 0 -1 2066
box -6 -6 124 52
use via__LI_M1  via__LI_M1_11
timestamp 1715010268
transform -1 0 807 0 -1 2066
box -6 -6 124 52
use via__LI_M1  via__LI_M1_12
timestamp 1715010268
transform -1 0 607 0 -1 2066
box -6 -6 124 52
use via__LI_M1  via__LI_M1_13
timestamp 1715010268
transform -1 0 407 0 -1 2066
box -6 -6 124 52
use via__LI_M1  via__LI_M1_14
timestamp 1715010268
transform 0 1 76 -1 0 1853
box -6 -6 124 52
use via__LI_M1  via__LI_M1_15
timestamp 1715010268
transform 0 1 76 -1 0 1653
box -6 -6 124 52
use via__LI_M1  via__LI_M1_16
timestamp 1715010268
transform 0 1 76 -1 0 1253
box -6 -6 124 52
use via__LI_M1  via__LI_M1_17
timestamp 1715010268
transform 0 1 76 -1 0 1453
box -6 -6 124 52
use via__LI_M1  via__LI_M1_18
timestamp 1715010268
transform 0 1 76 -1 0 1053
box -6 -6 124 52
use via__LI_M1  via__LI_M1_19
timestamp 1715010268
transform 1 0 331 0 1 70
box -6 -6 124 52
use via__LI_M1  via__LI_M1_20
timestamp 1715010268
transform 1 0 531 0 1 70
box -6 -6 124 52
use via__LI_M1  via__LI_M1_21
timestamp 1715010268
transform 1 0 731 0 1 70
box -6 -6 124 52
use via__LI_M1  via__LI_M1_22
timestamp 1715010268
transform 0 1 76 -1 0 653
box -6 -6 124 52
use via__LI_M1  via__LI_M1_23
timestamp 1715010268
transform 1 0 931 0 1 70
box -6 -6 124 52
use via__LI_M1  via__LI_M1_24
timestamp 1715010268
transform 1 0 1131 0 1 70
box -6 -6 124 52
use via__LI_M1  via__LI_M1_25
timestamp 1715010268
transform 0 1 76 -1 0 453
box -6 -6 124 52
use via__LI_M1  via__LI_M1_26
timestamp 1715010268
transform 0 1 76 -1 0 853
box -6 -6 124 52
use via__LI_M1  via__LI_M1_27
timestamp 1715010268
transform 0 -1 2476 1 0 990
box -6 -6 124 52
use via__LI_M1  via__LI_M1_28
timestamp 1715010268
transform 1 0 1331 0 1 70
box -6 -6 124 52
use via__LI_M1  via__LI_M1_29
timestamp 1715010268
transform 1 0 1531 0 1 70
box -6 -6 124 52
use via__LI_M1  via__LI_M1_30
timestamp 1715010268
transform 1 0 1731 0 1 70
box -6 -6 124 52
use via__LI_M1  via__LI_M1_31
timestamp 1715010268
transform 1 0 1931 0 1 70
box -6 -6 124 52
use via__LI_M1  via__LI_M1_32
timestamp 1715010268
transform 1 0 2131 0 1 70
box -6 -6 124 52
use via__LI_M1  via__LI_M1_33
timestamp 1715010268
transform 0 -1 2476 1 0 390
box -6 -6 124 52
use via__LI_M1  via__LI_M1_34
timestamp 1715010268
transform 0 -1 2476 1 0 590
box -6 -6 124 52
use via__LI_M1  via__LI_M1_35
timestamp 1715010268
transform 0 -1 2476 1 0 790
box -6 -6 124 52
use via__M1_M2  via__M1_M2_0
timestamp 1715010268
transform 0 -1 1582 1 0 833
box 0 0 140 80
use via__M1_M2  via__M1_M2_1
timestamp 1715010268
transform 0 -1 1066 1 0 833
box 0 0 140 80
use via__M1_M2  via__M1_M2_2
timestamp 1715010268
transform 0 -1 139 1 0 1141
box 0 0 140 80
use via__M1_M2  via__M1_M2_3
timestamp 1715010268
transform 0 -1 2256 1 0 1173
box 0 0 140 80
use via__M1_M2  via__M1_M2_4
timestamp 1715010268
transform 0 -1 139 1 0 1001
box 0 0 140 80
use via__M1_M2  via__M1_M2_5
timestamp 1715010268
transform 0 -1 139 1 0 861
box 0 0 140 80
use via__M1_M2  via__M1_M2_6
timestamp 1715010268
transform 0 -1 1740 1 0 1173
box 0 0 140 80
use via__M1_M2  via__M1_M2_7
timestamp 1715010268
transform 0 -1 1582 1 0 619
box 0 0 140 80
use via__M1_M2  via__M1_M2_8
timestamp 1715010268
transform 0 -1 1066 1 0 619
box 0 0 140 80
use via__M1_M2  via__M1_M2_9
timestamp 1715010268
transform 0 -1 908 1 0 1173
box 0 0 140 80
use via__M1_M2  via__M1_M2_10
timestamp 1715010268
transform 0 -1 392 1 0 1173
box 0 0 140 80
use via__M1_M2  via__M1_M2_11
timestamp 1715010268
transform 0 -1 1582 1 0 1387
box 0 0 140 80
use via__M1_M2  via__M1_M2_12
timestamp 1715010268
transform 0 -1 1066 1 0 1387
box 0 0 140 80
use via__M1_M2  via__M1_M2_13
timestamp 1715010268
transform 0 1 164 1 0 472
box 0 0 140 80
use via__M1_M2  via__M1_M2_14
timestamp 1715010268
transform 0 1 164 1 0 332
box 0 0 140 80
use via__M1_M2  via__M1_M2_15
timestamp 1715010268
transform 0 -1 1998 -1 0 1143
box 0 0 140 80
use via__M1_M2  via__M1_M2_16
timestamp 1715010268
transform 0 -1 1324 -1 0 1143
box 0 0 140 80
use via__M1_M2  via__M1_M2_17
timestamp 1715010268
transform 0 -1 650 -1 0 1143
box 0 0 140 80
use via__M2_M3  via__M2_M3_0
timestamp 1715010268
transform 0 1 986 -1 0 983
box 0 0 160 80
use via__M2_M3  via__M2_M3_1
timestamp 1715010268
transform 1 0 138 0 1 1032
box 0 0 160 80
use via__M2_M3  via__M2_M3_2
timestamp 1715010268
transform 0 1 1502 -1 0 983
box 0 0 160 80
<< labels >>
flabel metal2 s 2309 0 2389 40 1 FreeSans 200 0 0 0 vbn
port 3 nsew
flabel metal2 s 164 0 244 40 1 FreeSans 200 0 0 0 vbp
port 5 nsew
flabel metal3 s 2506 863 2549 943 1 FreeSans 200 0 0 0 ibp
port 8 nsew
flabel metal3 s 0 1032 46 1112 1 FreeSans 200 0 0 0 vdd
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 2549 2096
string path 2.475 26.800 49.200 26.800 
<< end >>
