magic
tech sky130A
magscale 1 2
timestamp 1715625863
<< pwell >>
rect -4085 1802 4085 1888
rect -4085 -1802 -3999 1802
rect 3999 -1802 4085 1802
rect -4085 -1888 4085 -1802
<< psubdiff >>
rect -4059 1828 -3961 1862
rect -3927 1828 -3893 1862
rect -3859 1828 -3825 1862
rect -3791 1828 -3757 1862
rect -3723 1828 -3689 1862
rect -3655 1828 -3621 1862
rect -3587 1828 -3553 1862
rect -3519 1828 -3485 1862
rect -3451 1828 -3417 1862
rect -3383 1828 -3349 1862
rect -3315 1828 -3281 1862
rect -3247 1828 -3213 1862
rect -3179 1828 -3145 1862
rect -3111 1828 -3077 1862
rect -3043 1828 -3009 1862
rect -2975 1828 -2941 1862
rect -2907 1828 -2873 1862
rect -2839 1828 -2805 1862
rect -2771 1828 -2737 1862
rect -2703 1828 -2669 1862
rect -2635 1828 -2601 1862
rect -2567 1828 -2533 1862
rect -2499 1828 -2465 1862
rect -2431 1828 -2397 1862
rect -2363 1828 -2329 1862
rect -2295 1828 -2261 1862
rect -2227 1828 -2193 1862
rect -2159 1828 -2125 1862
rect -2091 1828 -2057 1862
rect -2023 1828 -1989 1862
rect -1955 1828 -1921 1862
rect -1887 1828 -1853 1862
rect -1819 1828 -1785 1862
rect -1751 1828 -1717 1862
rect -1683 1828 -1649 1862
rect -1615 1828 -1581 1862
rect -1547 1828 -1513 1862
rect -1479 1828 -1445 1862
rect -1411 1828 -1377 1862
rect -1343 1828 -1309 1862
rect -1275 1828 -1241 1862
rect -1207 1828 -1173 1862
rect -1139 1828 -1105 1862
rect -1071 1828 -1037 1862
rect -1003 1828 -969 1862
rect -935 1828 -901 1862
rect -867 1828 -833 1862
rect -799 1828 -765 1862
rect -731 1828 -697 1862
rect -663 1828 -629 1862
rect -595 1828 -561 1862
rect -527 1828 -493 1862
rect -459 1828 -425 1862
rect -391 1828 -357 1862
rect -323 1828 -289 1862
rect -255 1828 -221 1862
rect -187 1828 -153 1862
rect -119 1828 -85 1862
rect -51 1828 -17 1862
rect 17 1828 51 1862
rect 85 1828 119 1862
rect 153 1828 187 1862
rect 221 1828 255 1862
rect 289 1828 323 1862
rect 357 1828 391 1862
rect 425 1828 459 1862
rect 493 1828 527 1862
rect 561 1828 595 1862
rect 629 1828 663 1862
rect 697 1828 731 1862
rect 765 1828 799 1862
rect 833 1828 867 1862
rect 901 1828 935 1862
rect 969 1828 1003 1862
rect 1037 1828 1071 1862
rect 1105 1828 1139 1862
rect 1173 1828 1207 1862
rect 1241 1828 1275 1862
rect 1309 1828 1343 1862
rect 1377 1828 1411 1862
rect 1445 1828 1479 1862
rect 1513 1828 1547 1862
rect 1581 1828 1615 1862
rect 1649 1828 1683 1862
rect 1717 1828 1751 1862
rect 1785 1828 1819 1862
rect 1853 1828 1887 1862
rect 1921 1828 1955 1862
rect 1989 1828 2023 1862
rect 2057 1828 2091 1862
rect 2125 1828 2159 1862
rect 2193 1828 2227 1862
rect 2261 1828 2295 1862
rect 2329 1828 2363 1862
rect 2397 1828 2431 1862
rect 2465 1828 2499 1862
rect 2533 1828 2567 1862
rect 2601 1828 2635 1862
rect 2669 1828 2703 1862
rect 2737 1828 2771 1862
rect 2805 1828 2839 1862
rect 2873 1828 2907 1862
rect 2941 1828 2975 1862
rect 3009 1828 3043 1862
rect 3077 1828 3111 1862
rect 3145 1828 3179 1862
rect 3213 1828 3247 1862
rect 3281 1828 3315 1862
rect 3349 1828 3383 1862
rect 3417 1828 3451 1862
rect 3485 1828 3519 1862
rect 3553 1828 3587 1862
rect 3621 1828 3655 1862
rect 3689 1828 3723 1862
rect 3757 1828 3791 1862
rect 3825 1828 3859 1862
rect 3893 1828 3927 1862
rect 3961 1828 4059 1862
rect -4059 1751 -4025 1828
rect 4025 1751 4059 1828
rect -4059 1683 -4025 1717
rect -4059 1615 -4025 1649
rect -4059 1547 -4025 1581
rect -4059 1479 -4025 1513
rect -4059 1411 -4025 1445
rect -4059 1343 -4025 1377
rect -4059 1275 -4025 1309
rect -4059 1207 -4025 1241
rect -4059 1139 -4025 1173
rect -4059 1071 -4025 1105
rect -4059 1003 -4025 1037
rect -4059 935 -4025 969
rect -4059 867 -4025 901
rect -4059 799 -4025 833
rect -4059 731 -4025 765
rect -4059 663 -4025 697
rect -4059 595 -4025 629
rect -4059 527 -4025 561
rect -4059 459 -4025 493
rect -4059 391 -4025 425
rect -4059 323 -4025 357
rect -4059 255 -4025 289
rect -4059 187 -4025 221
rect -4059 119 -4025 153
rect -4059 51 -4025 85
rect -4059 -17 -4025 17
rect -4059 -85 -4025 -51
rect -4059 -153 -4025 -119
rect -4059 -221 -4025 -187
rect -4059 -289 -4025 -255
rect -4059 -357 -4025 -323
rect -4059 -425 -4025 -391
rect -4059 -493 -4025 -459
rect -4059 -561 -4025 -527
rect -4059 -629 -4025 -595
rect -4059 -697 -4025 -663
rect -4059 -765 -4025 -731
rect -4059 -833 -4025 -799
rect -4059 -901 -4025 -867
rect -4059 -969 -4025 -935
rect -4059 -1037 -4025 -1003
rect -4059 -1105 -4025 -1071
rect -4059 -1173 -4025 -1139
rect -4059 -1241 -4025 -1207
rect -4059 -1309 -4025 -1275
rect -4059 -1377 -4025 -1343
rect -4059 -1445 -4025 -1411
rect -4059 -1513 -4025 -1479
rect -4059 -1581 -4025 -1547
rect -4059 -1649 -4025 -1615
rect -4059 -1717 -4025 -1683
rect 4025 1683 4059 1717
rect 4025 1615 4059 1649
rect 4025 1547 4059 1581
rect 4025 1479 4059 1513
rect 4025 1411 4059 1445
rect 4025 1343 4059 1377
rect 4025 1275 4059 1309
rect 4025 1207 4059 1241
rect 4025 1139 4059 1173
rect 4025 1071 4059 1105
rect 4025 1003 4059 1037
rect 4025 935 4059 969
rect 4025 867 4059 901
rect 4025 799 4059 833
rect 4025 731 4059 765
rect 4025 663 4059 697
rect 4025 595 4059 629
rect 4025 527 4059 561
rect 4025 459 4059 493
rect 4025 391 4059 425
rect 4025 323 4059 357
rect 4025 255 4059 289
rect 4025 187 4059 221
rect 4025 119 4059 153
rect 4025 51 4059 85
rect 4025 -17 4059 17
rect 4025 -85 4059 -51
rect 4025 -153 4059 -119
rect 4025 -221 4059 -187
rect 4025 -289 4059 -255
rect 4025 -357 4059 -323
rect 4025 -425 4059 -391
rect 4025 -493 4059 -459
rect 4025 -561 4059 -527
rect 4025 -629 4059 -595
rect 4025 -697 4059 -663
rect 4025 -765 4059 -731
rect 4025 -833 4059 -799
rect 4025 -901 4059 -867
rect 4025 -969 4059 -935
rect 4025 -1037 4059 -1003
rect 4025 -1105 4059 -1071
rect 4025 -1173 4059 -1139
rect 4025 -1241 4059 -1207
rect 4025 -1309 4059 -1275
rect 4025 -1377 4059 -1343
rect 4025 -1445 4059 -1411
rect 4025 -1513 4059 -1479
rect 4025 -1581 4059 -1547
rect 4025 -1649 4059 -1615
rect 4025 -1717 4059 -1683
rect -4059 -1828 -4025 -1751
rect 4025 -1828 4059 -1751
rect -4059 -1862 -3961 -1828
rect -3927 -1862 -3893 -1828
rect -3859 -1862 -3825 -1828
rect -3791 -1862 -3757 -1828
rect -3723 -1862 -3689 -1828
rect -3655 -1862 -3621 -1828
rect -3587 -1862 -3553 -1828
rect -3519 -1862 -3485 -1828
rect -3451 -1862 -3417 -1828
rect -3383 -1862 -3349 -1828
rect -3315 -1862 -3281 -1828
rect -3247 -1862 -3213 -1828
rect -3179 -1862 -3145 -1828
rect -3111 -1862 -3077 -1828
rect -3043 -1862 -3009 -1828
rect -2975 -1862 -2941 -1828
rect -2907 -1862 -2873 -1828
rect -2839 -1862 -2805 -1828
rect -2771 -1862 -2737 -1828
rect -2703 -1862 -2669 -1828
rect -2635 -1862 -2601 -1828
rect -2567 -1862 -2533 -1828
rect -2499 -1862 -2465 -1828
rect -2431 -1862 -2397 -1828
rect -2363 -1862 -2329 -1828
rect -2295 -1862 -2261 -1828
rect -2227 -1862 -2193 -1828
rect -2159 -1862 -2125 -1828
rect -2091 -1862 -2057 -1828
rect -2023 -1862 -1989 -1828
rect -1955 -1862 -1921 -1828
rect -1887 -1862 -1853 -1828
rect -1819 -1862 -1785 -1828
rect -1751 -1862 -1717 -1828
rect -1683 -1862 -1649 -1828
rect -1615 -1862 -1581 -1828
rect -1547 -1862 -1513 -1828
rect -1479 -1862 -1445 -1828
rect -1411 -1862 -1377 -1828
rect -1343 -1862 -1309 -1828
rect -1275 -1862 -1241 -1828
rect -1207 -1862 -1173 -1828
rect -1139 -1862 -1105 -1828
rect -1071 -1862 -1037 -1828
rect -1003 -1862 -969 -1828
rect -935 -1862 -901 -1828
rect -867 -1862 -833 -1828
rect -799 -1862 -765 -1828
rect -731 -1862 -697 -1828
rect -663 -1862 -629 -1828
rect -595 -1862 -561 -1828
rect -527 -1862 -493 -1828
rect -459 -1862 -425 -1828
rect -391 -1862 -357 -1828
rect -323 -1862 -289 -1828
rect -255 -1862 -221 -1828
rect -187 -1862 -153 -1828
rect -119 -1862 -85 -1828
rect -51 -1862 -17 -1828
rect 17 -1862 51 -1828
rect 85 -1862 119 -1828
rect 153 -1862 187 -1828
rect 221 -1862 255 -1828
rect 289 -1862 323 -1828
rect 357 -1862 391 -1828
rect 425 -1862 459 -1828
rect 493 -1862 527 -1828
rect 561 -1862 595 -1828
rect 629 -1862 663 -1828
rect 697 -1862 731 -1828
rect 765 -1862 799 -1828
rect 833 -1862 867 -1828
rect 901 -1862 935 -1828
rect 969 -1862 1003 -1828
rect 1037 -1862 1071 -1828
rect 1105 -1862 1139 -1828
rect 1173 -1862 1207 -1828
rect 1241 -1862 1275 -1828
rect 1309 -1862 1343 -1828
rect 1377 -1862 1411 -1828
rect 1445 -1862 1479 -1828
rect 1513 -1862 1547 -1828
rect 1581 -1862 1615 -1828
rect 1649 -1862 1683 -1828
rect 1717 -1862 1751 -1828
rect 1785 -1862 1819 -1828
rect 1853 -1862 1887 -1828
rect 1921 -1862 1955 -1828
rect 1989 -1862 2023 -1828
rect 2057 -1862 2091 -1828
rect 2125 -1862 2159 -1828
rect 2193 -1862 2227 -1828
rect 2261 -1862 2295 -1828
rect 2329 -1862 2363 -1828
rect 2397 -1862 2431 -1828
rect 2465 -1862 2499 -1828
rect 2533 -1862 2567 -1828
rect 2601 -1862 2635 -1828
rect 2669 -1862 2703 -1828
rect 2737 -1862 2771 -1828
rect 2805 -1862 2839 -1828
rect 2873 -1862 2907 -1828
rect 2941 -1862 2975 -1828
rect 3009 -1862 3043 -1828
rect 3077 -1862 3111 -1828
rect 3145 -1862 3179 -1828
rect 3213 -1862 3247 -1828
rect 3281 -1862 3315 -1828
rect 3349 -1862 3383 -1828
rect 3417 -1862 3451 -1828
rect 3485 -1862 3519 -1828
rect 3553 -1862 3587 -1828
rect 3621 -1862 3655 -1828
rect 3689 -1862 3723 -1828
rect 3757 -1862 3791 -1828
rect 3825 -1862 3859 -1828
rect 3893 -1862 3927 -1828
rect 3961 -1862 4059 -1828
<< psubdiffcont >>
rect -3961 1828 -3927 1862
rect -3893 1828 -3859 1862
rect -3825 1828 -3791 1862
rect -3757 1828 -3723 1862
rect -3689 1828 -3655 1862
rect -3621 1828 -3587 1862
rect -3553 1828 -3519 1862
rect -3485 1828 -3451 1862
rect -3417 1828 -3383 1862
rect -3349 1828 -3315 1862
rect -3281 1828 -3247 1862
rect -3213 1828 -3179 1862
rect -3145 1828 -3111 1862
rect -3077 1828 -3043 1862
rect -3009 1828 -2975 1862
rect -2941 1828 -2907 1862
rect -2873 1828 -2839 1862
rect -2805 1828 -2771 1862
rect -2737 1828 -2703 1862
rect -2669 1828 -2635 1862
rect -2601 1828 -2567 1862
rect -2533 1828 -2499 1862
rect -2465 1828 -2431 1862
rect -2397 1828 -2363 1862
rect -2329 1828 -2295 1862
rect -2261 1828 -2227 1862
rect -2193 1828 -2159 1862
rect -2125 1828 -2091 1862
rect -2057 1828 -2023 1862
rect -1989 1828 -1955 1862
rect -1921 1828 -1887 1862
rect -1853 1828 -1819 1862
rect -1785 1828 -1751 1862
rect -1717 1828 -1683 1862
rect -1649 1828 -1615 1862
rect -1581 1828 -1547 1862
rect -1513 1828 -1479 1862
rect -1445 1828 -1411 1862
rect -1377 1828 -1343 1862
rect -1309 1828 -1275 1862
rect -1241 1828 -1207 1862
rect -1173 1828 -1139 1862
rect -1105 1828 -1071 1862
rect -1037 1828 -1003 1862
rect -969 1828 -935 1862
rect -901 1828 -867 1862
rect -833 1828 -799 1862
rect -765 1828 -731 1862
rect -697 1828 -663 1862
rect -629 1828 -595 1862
rect -561 1828 -527 1862
rect -493 1828 -459 1862
rect -425 1828 -391 1862
rect -357 1828 -323 1862
rect -289 1828 -255 1862
rect -221 1828 -187 1862
rect -153 1828 -119 1862
rect -85 1828 -51 1862
rect -17 1828 17 1862
rect 51 1828 85 1862
rect 119 1828 153 1862
rect 187 1828 221 1862
rect 255 1828 289 1862
rect 323 1828 357 1862
rect 391 1828 425 1862
rect 459 1828 493 1862
rect 527 1828 561 1862
rect 595 1828 629 1862
rect 663 1828 697 1862
rect 731 1828 765 1862
rect 799 1828 833 1862
rect 867 1828 901 1862
rect 935 1828 969 1862
rect 1003 1828 1037 1862
rect 1071 1828 1105 1862
rect 1139 1828 1173 1862
rect 1207 1828 1241 1862
rect 1275 1828 1309 1862
rect 1343 1828 1377 1862
rect 1411 1828 1445 1862
rect 1479 1828 1513 1862
rect 1547 1828 1581 1862
rect 1615 1828 1649 1862
rect 1683 1828 1717 1862
rect 1751 1828 1785 1862
rect 1819 1828 1853 1862
rect 1887 1828 1921 1862
rect 1955 1828 1989 1862
rect 2023 1828 2057 1862
rect 2091 1828 2125 1862
rect 2159 1828 2193 1862
rect 2227 1828 2261 1862
rect 2295 1828 2329 1862
rect 2363 1828 2397 1862
rect 2431 1828 2465 1862
rect 2499 1828 2533 1862
rect 2567 1828 2601 1862
rect 2635 1828 2669 1862
rect 2703 1828 2737 1862
rect 2771 1828 2805 1862
rect 2839 1828 2873 1862
rect 2907 1828 2941 1862
rect 2975 1828 3009 1862
rect 3043 1828 3077 1862
rect 3111 1828 3145 1862
rect 3179 1828 3213 1862
rect 3247 1828 3281 1862
rect 3315 1828 3349 1862
rect 3383 1828 3417 1862
rect 3451 1828 3485 1862
rect 3519 1828 3553 1862
rect 3587 1828 3621 1862
rect 3655 1828 3689 1862
rect 3723 1828 3757 1862
rect 3791 1828 3825 1862
rect 3859 1828 3893 1862
rect 3927 1828 3961 1862
rect -4059 1717 -4025 1751
rect -4059 1649 -4025 1683
rect -4059 1581 -4025 1615
rect -4059 1513 -4025 1547
rect -4059 1445 -4025 1479
rect -4059 1377 -4025 1411
rect -4059 1309 -4025 1343
rect -4059 1241 -4025 1275
rect -4059 1173 -4025 1207
rect -4059 1105 -4025 1139
rect -4059 1037 -4025 1071
rect -4059 969 -4025 1003
rect -4059 901 -4025 935
rect -4059 833 -4025 867
rect -4059 765 -4025 799
rect -4059 697 -4025 731
rect -4059 629 -4025 663
rect -4059 561 -4025 595
rect -4059 493 -4025 527
rect -4059 425 -4025 459
rect -4059 357 -4025 391
rect -4059 289 -4025 323
rect -4059 221 -4025 255
rect -4059 153 -4025 187
rect -4059 85 -4025 119
rect -4059 17 -4025 51
rect -4059 -51 -4025 -17
rect -4059 -119 -4025 -85
rect -4059 -187 -4025 -153
rect -4059 -255 -4025 -221
rect -4059 -323 -4025 -289
rect -4059 -391 -4025 -357
rect -4059 -459 -4025 -425
rect -4059 -527 -4025 -493
rect -4059 -595 -4025 -561
rect -4059 -663 -4025 -629
rect -4059 -731 -4025 -697
rect -4059 -799 -4025 -765
rect -4059 -867 -4025 -833
rect -4059 -935 -4025 -901
rect -4059 -1003 -4025 -969
rect -4059 -1071 -4025 -1037
rect -4059 -1139 -4025 -1105
rect -4059 -1207 -4025 -1173
rect -4059 -1275 -4025 -1241
rect -4059 -1343 -4025 -1309
rect -4059 -1411 -4025 -1377
rect -4059 -1479 -4025 -1445
rect -4059 -1547 -4025 -1513
rect -4059 -1615 -4025 -1581
rect -4059 -1683 -4025 -1649
rect -4059 -1751 -4025 -1717
rect 4025 1717 4059 1751
rect 4025 1649 4059 1683
rect 4025 1581 4059 1615
rect 4025 1513 4059 1547
rect 4025 1445 4059 1479
rect 4025 1377 4059 1411
rect 4025 1309 4059 1343
rect 4025 1241 4059 1275
rect 4025 1173 4059 1207
rect 4025 1105 4059 1139
rect 4025 1037 4059 1071
rect 4025 969 4059 1003
rect 4025 901 4059 935
rect 4025 833 4059 867
rect 4025 765 4059 799
rect 4025 697 4059 731
rect 4025 629 4059 663
rect 4025 561 4059 595
rect 4025 493 4059 527
rect 4025 425 4059 459
rect 4025 357 4059 391
rect 4025 289 4059 323
rect 4025 221 4059 255
rect 4025 153 4059 187
rect 4025 85 4059 119
rect 4025 17 4059 51
rect 4025 -51 4059 -17
rect 4025 -119 4059 -85
rect 4025 -187 4059 -153
rect 4025 -255 4059 -221
rect 4025 -323 4059 -289
rect 4025 -391 4059 -357
rect 4025 -459 4059 -425
rect 4025 -527 4059 -493
rect 4025 -595 4059 -561
rect 4025 -663 4059 -629
rect 4025 -731 4059 -697
rect 4025 -799 4059 -765
rect 4025 -867 4059 -833
rect 4025 -935 4059 -901
rect 4025 -1003 4059 -969
rect 4025 -1071 4059 -1037
rect 4025 -1139 4059 -1105
rect 4025 -1207 4059 -1173
rect 4025 -1275 4059 -1241
rect 4025 -1343 4059 -1309
rect 4025 -1411 4059 -1377
rect 4025 -1479 4059 -1445
rect 4025 -1547 4059 -1513
rect 4025 -1615 4059 -1581
rect 4025 -1683 4059 -1649
rect 4025 -1751 4059 -1717
rect -3961 -1862 -3927 -1828
rect -3893 -1862 -3859 -1828
rect -3825 -1862 -3791 -1828
rect -3757 -1862 -3723 -1828
rect -3689 -1862 -3655 -1828
rect -3621 -1862 -3587 -1828
rect -3553 -1862 -3519 -1828
rect -3485 -1862 -3451 -1828
rect -3417 -1862 -3383 -1828
rect -3349 -1862 -3315 -1828
rect -3281 -1862 -3247 -1828
rect -3213 -1862 -3179 -1828
rect -3145 -1862 -3111 -1828
rect -3077 -1862 -3043 -1828
rect -3009 -1862 -2975 -1828
rect -2941 -1862 -2907 -1828
rect -2873 -1862 -2839 -1828
rect -2805 -1862 -2771 -1828
rect -2737 -1862 -2703 -1828
rect -2669 -1862 -2635 -1828
rect -2601 -1862 -2567 -1828
rect -2533 -1862 -2499 -1828
rect -2465 -1862 -2431 -1828
rect -2397 -1862 -2363 -1828
rect -2329 -1862 -2295 -1828
rect -2261 -1862 -2227 -1828
rect -2193 -1862 -2159 -1828
rect -2125 -1862 -2091 -1828
rect -2057 -1862 -2023 -1828
rect -1989 -1862 -1955 -1828
rect -1921 -1862 -1887 -1828
rect -1853 -1862 -1819 -1828
rect -1785 -1862 -1751 -1828
rect -1717 -1862 -1683 -1828
rect -1649 -1862 -1615 -1828
rect -1581 -1862 -1547 -1828
rect -1513 -1862 -1479 -1828
rect -1445 -1862 -1411 -1828
rect -1377 -1862 -1343 -1828
rect -1309 -1862 -1275 -1828
rect -1241 -1862 -1207 -1828
rect -1173 -1862 -1139 -1828
rect -1105 -1862 -1071 -1828
rect -1037 -1862 -1003 -1828
rect -969 -1862 -935 -1828
rect -901 -1862 -867 -1828
rect -833 -1862 -799 -1828
rect -765 -1862 -731 -1828
rect -697 -1862 -663 -1828
rect -629 -1862 -595 -1828
rect -561 -1862 -527 -1828
rect -493 -1862 -459 -1828
rect -425 -1862 -391 -1828
rect -357 -1862 -323 -1828
rect -289 -1862 -255 -1828
rect -221 -1862 -187 -1828
rect -153 -1862 -119 -1828
rect -85 -1862 -51 -1828
rect -17 -1862 17 -1828
rect 51 -1862 85 -1828
rect 119 -1862 153 -1828
rect 187 -1862 221 -1828
rect 255 -1862 289 -1828
rect 323 -1862 357 -1828
rect 391 -1862 425 -1828
rect 459 -1862 493 -1828
rect 527 -1862 561 -1828
rect 595 -1862 629 -1828
rect 663 -1862 697 -1828
rect 731 -1862 765 -1828
rect 799 -1862 833 -1828
rect 867 -1862 901 -1828
rect 935 -1862 969 -1828
rect 1003 -1862 1037 -1828
rect 1071 -1862 1105 -1828
rect 1139 -1862 1173 -1828
rect 1207 -1862 1241 -1828
rect 1275 -1862 1309 -1828
rect 1343 -1862 1377 -1828
rect 1411 -1862 1445 -1828
rect 1479 -1862 1513 -1828
rect 1547 -1862 1581 -1828
rect 1615 -1862 1649 -1828
rect 1683 -1862 1717 -1828
rect 1751 -1862 1785 -1828
rect 1819 -1862 1853 -1828
rect 1887 -1862 1921 -1828
rect 1955 -1862 1989 -1828
rect 2023 -1862 2057 -1828
rect 2091 -1862 2125 -1828
rect 2159 -1862 2193 -1828
rect 2227 -1862 2261 -1828
rect 2295 -1862 2329 -1828
rect 2363 -1862 2397 -1828
rect 2431 -1862 2465 -1828
rect 2499 -1862 2533 -1828
rect 2567 -1862 2601 -1828
rect 2635 -1862 2669 -1828
rect 2703 -1862 2737 -1828
rect 2771 -1862 2805 -1828
rect 2839 -1862 2873 -1828
rect 2907 -1862 2941 -1828
rect 2975 -1862 3009 -1828
rect 3043 -1862 3077 -1828
rect 3111 -1862 3145 -1828
rect 3179 -1862 3213 -1828
rect 3247 -1862 3281 -1828
rect 3315 -1862 3349 -1828
rect 3383 -1862 3417 -1828
rect 3451 -1862 3485 -1828
rect 3519 -1862 3553 -1828
rect 3587 -1862 3621 -1828
rect 3655 -1862 3689 -1828
rect 3723 -1862 3757 -1828
rect 3791 -1862 3825 -1828
rect 3859 -1862 3893 -1828
rect 3927 -1862 3961 -1828
<< xpolycontact >>
rect -3929 1296 -3791 1732
rect -3929 -1732 -3791 -1296
rect -3543 1296 -3405 1732
rect -3543 -1732 -3405 -1296
rect -3157 1296 -3019 1732
rect -3157 -1732 -3019 -1296
rect -2771 1296 -2633 1732
rect -2771 -1732 -2633 -1296
rect -2385 1296 -2247 1732
rect -2385 -1732 -2247 -1296
rect -1999 1296 -1861 1732
rect -1999 -1732 -1861 -1296
rect -1613 1296 -1475 1732
rect -1613 -1732 -1475 -1296
rect -1227 1296 -1089 1732
rect -1227 -1732 -1089 -1296
rect -841 1296 -703 1732
rect -841 -1732 -703 -1296
rect -455 1296 -317 1732
rect -455 -1732 -317 -1296
rect -69 1296 69 1732
rect -69 -1732 69 -1296
rect 317 1296 455 1732
rect 317 -1732 455 -1296
rect 703 1296 841 1732
rect 703 -1732 841 -1296
rect 1089 1296 1227 1732
rect 1089 -1732 1227 -1296
rect 1475 1296 1613 1732
rect 1475 -1732 1613 -1296
rect 1861 1296 1999 1732
rect 1861 -1732 1999 -1296
rect 2247 1296 2385 1732
rect 2247 -1732 2385 -1296
rect 2633 1296 2771 1732
rect 2633 -1732 2771 -1296
rect 3019 1296 3157 1732
rect 3019 -1732 3157 -1296
rect 3405 1296 3543 1732
rect 3405 -1732 3543 -1296
rect 3791 1296 3929 1732
rect 3791 -1732 3929 -1296
<< xpolyres >>
rect -3929 -1296 -3791 1296
rect -3543 -1296 -3405 1296
rect -3157 -1296 -3019 1296
rect -2771 -1296 -2633 1296
rect -2385 -1296 -2247 1296
rect -1999 -1296 -1861 1296
rect -1613 -1296 -1475 1296
rect -1227 -1296 -1089 1296
rect -841 -1296 -703 1296
rect -455 -1296 -317 1296
rect -69 -1296 69 1296
rect 317 -1296 455 1296
rect 703 -1296 841 1296
rect 1089 -1296 1227 1296
rect 1475 -1296 1613 1296
rect 1861 -1296 1999 1296
rect 2247 -1296 2385 1296
rect 2633 -1296 2771 1296
rect 3019 -1296 3157 1296
rect 3405 -1296 3543 1296
rect 3791 -1296 3929 1296
<< locali >>
rect -4059 1828 -3961 1862
rect -3927 1828 -3893 1862
rect -3859 1828 -3825 1862
rect -3791 1828 -3757 1862
rect -3723 1828 -3689 1862
rect -3655 1828 -3621 1862
rect -3587 1828 -3553 1862
rect -3519 1828 -3485 1862
rect -3451 1828 -3417 1862
rect -3383 1828 -3349 1862
rect -3315 1828 -3281 1862
rect -3247 1828 -3213 1862
rect -3179 1828 -3145 1862
rect -3111 1828 -3077 1862
rect -3043 1828 -3009 1862
rect -2975 1828 -2941 1862
rect -2907 1828 -2873 1862
rect -2839 1828 -2805 1862
rect -2771 1828 -2737 1862
rect -2703 1828 -2669 1862
rect -2635 1828 -2601 1862
rect -2567 1828 -2533 1862
rect -2499 1828 -2465 1862
rect -2431 1828 -2397 1862
rect -2363 1828 -2329 1862
rect -2295 1828 -2261 1862
rect -2227 1828 -2193 1862
rect -2159 1828 -2125 1862
rect -2091 1828 -2057 1862
rect -2023 1828 -1989 1862
rect -1955 1828 -1921 1862
rect -1887 1828 -1853 1862
rect -1819 1828 -1785 1862
rect -1751 1828 -1717 1862
rect -1683 1828 -1649 1862
rect -1615 1828 -1581 1862
rect -1547 1828 -1513 1862
rect -1479 1828 -1445 1862
rect -1411 1828 -1377 1862
rect -1343 1828 -1309 1862
rect -1275 1828 -1241 1862
rect -1207 1828 -1173 1862
rect -1139 1828 -1105 1862
rect -1071 1828 -1037 1862
rect -1003 1828 -969 1862
rect -935 1828 -901 1862
rect -867 1828 -833 1862
rect -799 1828 -765 1862
rect -731 1828 -697 1862
rect -663 1828 -629 1862
rect -595 1828 -561 1862
rect -527 1828 -493 1862
rect -459 1828 -425 1862
rect -391 1828 -357 1862
rect -323 1828 -289 1862
rect -255 1828 -221 1862
rect -187 1828 -153 1862
rect -119 1828 -85 1862
rect -51 1828 -17 1862
rect 17 1828 51 1862
rect 85 1828 119 1862
rect 153 1828 187 1862
rect 221 1828 255 1862
rect 289 1828 323 1862
rect 357 1828 391 1862
rect 425 1828 459 1862
rect 493 1828 527 1862
rect 561 1828 595 1862
rect 629 1828 663 1862
rect 697 1828 731 1862
rect 765 1828 799 1862
rect 833 1828 867 1862
rect 901 1828 935 1862
rect 969 1828 1003 1862
rect 1037 1828 1071 1862
rect 1105 1828 1139 1862
rect 1173 1828 1207 1862
rect 1241 1828 1275 1862
rect 1309 1828 1343 1862
rect 1377 1828 1411 1862
rect 1445 1828 1479 1862
rect 1513 1828 1547 1862
rect 1581 1828 1615 1862
rect 1649 1828 1683 1862
rect 1717 1828 1751 1862
rect 1785 1828 1819 1862
rect 1853 1828 1887 1862
rect 1921 1828 1955 1862
rect 1989 1828 2023 1862
rect 2057 1828 2091 1862
rect 2125 1828 2159 1862
rect 2193 1828 2227 1862
rect 2261 1828 2295 1862
rect 2329 1828 2363 1862
rect 2397 1828 2431 1862
rect 2465 1828 2499 1862
rect 2533 1828 2567 1862
rect 2601 1828 2635 1862
rect 2669 1828 2703 1862
rect 2737 1828 2771 1862
rect 2805 1828 2839 1862
rect 2873 1828 2907 1862
rect 2941 1828 2975 1862
rect 3009 1828 3043 1862
rect 3077 1828 3111 1862
rect 3145 1828 3179 1862
rect 3213 1828 3247 1862
rect 3281 1828 3315 1862
rect 3349 1828 3383 1862
rect 3417 1828 3451 1862
rect 3485 1828 3519 1862
rect 3553 1828 3587 1862
rect 3621 1828 3655 1862
rect 3689 1828 3723 1862
rect 3757 1828 3791 1862
rect 3825 1828 3859 1862
rect 3893 1828 3927 1862
rect 3961 1828 4059 1862
rect -4059 1751 -4025 1828
rect 4025 1751 4059 1828
rect -4059 1683 -4025 1717
rect -4059 1615 -4025 1649
rect -4059 1547 -4025 1581
rect -4059 1479 -4025 1513
rect -4059 1411 -4025 1445
rect -4059 1343 -4025 1377
rect -4059 1275 -4025 1309
rect 4025 1683 4059 1717
rect 4025 1615 4059 1649
rect 4025 1547 4059 1581
rect 4025 1479 4059 1513
rect 4025 1411 4059 1445
rect 4025 1343 4059 1377
rect -4059 1207 -4025 1241
rect -4059 1139 -4025 1173
rect -4059 1071 -4025 1105
rect -4059 1003 -4025 1037
rect -4059 935 -4025 969
rect -4059 867 -4025 901
rect -4059 799 -4025 833
rect -4059 731 -4025 765
rect -4059 663 -4025 697
rect -4059 595 -4025 629
rect -4059 527 -4025 561
rect -4059 459 -4025 493
rect -4059 391 -4025 425
rect -4059 323 -4025 357
rect -4059 255 -4025 289
rect -4059 187 -4025 221
rect -4059 119 -4025 153
rect -4059 51 -4025 85
rect -4059 -17 -4025 17
rect -4059 -85 -4025 -51
rect -4059 -153 -4025 -119
rect -4059 -221 -4025 -187
rect -4059 -289 -4025 -255
rect -4059 -357 -4025 -323
rect -4059 -425 -4025 -391
rect -4059 -493 -4025 -459
rect -4059 -561 -4025 -527
rect -4059 -629 -4025 -595
rect -4059 -697 -4025 -663
rect -4059 -765 -4025 -731
rect -4059 -833 -4025 -799
rect -4059 -901 -4025 -867
rect -4059 -969 -4025 -935
rect -4059 -1037 -4025 -1003
rect -4059 -1105 -4025 -1071
rect -4059 -1173 -4025 -1139
rect -4059 -1241 -4025 -1207
rect -4059 -1309 -4025 -1275
rect 4025 1275 4059 1309
rect 4025 1207 4059 1241
rect 4025 1139 4059 1173
rect 4025 1071 4059 1105
rect 4025 1003 4059 1037
rect 4025 935 4059 969
rect 4025 867 4059 901
rect 4025 799 4059 833
rect 4025 731 4059 765
rect 4025 663 4059 697
rect 4025 595 4059 629
rect 4025 527 4059 561
rect 4025 459 4059 493
rect 4025 391 4059 425
rect 4025 323 4059 357
rect 4025 255 4059 289
rect 4025 187 4059 221
rect 4025 119 4059 153
rect 4025 51 4059 85
rect 4025 -17 4059 17
rect 4025 -85 4059 -51
rect 4025 -153 4059 -119
rect 4025 -221 4059 -187
rect 4025 -289 4059 -255
rect 4025 -357 4059 -323
rect 4025 -425 4059 -391
rect 4025 -493 4059 -459
rect 4025 -561 4059 -527
rect 4025 -629 4059 -595
rect 4025 -697 4059 -663
rect 4025 -765 4059 -731
rect 4025 -833 4059 -799
rect 4025 -901 4059 -867
rect 4025 -969 4059 -935
rect 4025 -1037 4059 -1003
rect 4025 -1105 4059 -1071
rect 4025 -1173 4059 -1139
rect 4025 -1241 4059 -1207
rect -4059 -1377 -4025 -1343
rect -4059 -1445 -4025 -1411
rect -4059 -1513 -4025 -1479
rect -4059 -1581 -4025 -1547
rect -4059 -1649 -4025 -1615
rect -4059 -1717 -4025 -1683
rect 4025 -1309 4059 -1275
rect 4025 -1377 4059 -1343
rect 4025 -1445 4059 -1411
rect 4025 -1513 4059 -1479
rect 4025 -1581 4059 -1547
rect 4025 -1649 4059 -1615
rect 4025 -1717 4059 -1683
rect -4059 -1828 -4025 -1751
rect 4025 -1828 4059 -1751
rect -4059 -1862 -3961 -1828
rect -3927 -1862 -3893 -1828
rect -3859 -1862 -3825 -1828
rect -3791 -1862 -3757 -1828
rect -3723 -1862 -3689 -1828
rect -3655 -1862 -3621 -1828
rect -3587 -1862 -3553 -1828
rect -3519 -1862 -3485 -1828
rect -3451 -1862 -3417 -1828
rect -3383 -1862 -3349 -1828
rect -3315 -1862 -3281 -1828
rect -3247 -1862 -3213 -1828
rect -3179 -1862 -3145 -1828
rect -3111 -1862 -3077 -1828
rect -3043 -1862 -3009 -1828
rect -2975 -1862 -2941 -1828
rect -2907 -1862 -2873 -1828
rect -2839 -1862 -2805 -1828
rect -2771 -1862 -2737 -1828
rect -2703 -1862 -2669 -1828
rect -2635 -1862 -2601 -1828
rect -2567 -1862 -2533 -1828
rect -2499 -1862 -2465 -1828
rect -2431 -1862 -2397 -1828
rect -2363 -1862 -2329 -1828
rect -2295 -1862 -2261 -1828
rect -2227 -1862 -2193 -1828
rect -2159 -1862 -2125 -1828
rect -2091 -1862 -2057 -1828
rect -2023 -1862 -1989 -1828
rect -1955 -1862 -1921 -1828
rect -1887 -1862 -1853 -1828
rect -1819 -1862 -1785 -1828
rect -1751 -1862 -1717 -1828
rect -1683 -1862 -1649 -1828
rect -1615 -1862 -1581 -1828
rect -1547 -1862 -1513 -1828
rect -1479 -1862 -1445 -1828
rect -1411 -1862 -1377 -1828
rect -1343 -1862 -1309 -1828
rect -1275 -1862 -1241 -1828
rect -1207 -1862 -1173 -1828
rect -1139 -1862 -1105 -1828
rect -1071 -1862 -1037 -1828
rect -1003 -1862 -969 -1828
rect -935 -1862 -901 -1828
rect -867 -1862 -833 -1828
rect -799 -1862 -765 -1828
rect -731 -1862 -697 -1828
rect -663 -1862 -629 -1828
rect -595 -1862 -561 -1828
rect -527 -1862 -493 -1828
rect -459 -1862 -425 -1828
rect -391 -1862 -357 -1828
rect -323 -1862 -289 -1828
rect -255 -1862 -221 -1828
rect -187 -1862 -153 -1828
rect -119 -1862 -85 -1828
rect -51 -1862 -17 -1828
rect 17 -1862 51 -1828
rect 85 -1862 119 -1828
rect 153 -1862 187 -1828
rect 221 -1862 255 -1828
rect 289 -1862 323 -1828
rect 357 -1862 391 -1828
rect 425 -1862 459 -1828
rect 493 -1862 527 -1828
rect 561 -1862 595 -1828
rect 629 -1862 663 -1828
rect 697 -1862 731 -1828
rect 765 -1862 799 -1828
rect 833 -1862 867 -1828
rect 901 -1862 935 -1828
rect 969 -1862 1003 -1828
rect 1037 -1862 1071 -1828
rect 1105 -1862 1139 -1828
rect 1173 -1862 1207 -1828
rect 1241 -1862 1275 -1828
rect 1309 -1862 1343 -1828
rect 1377 -1862 1411 -1828
rect 1445 -1862 1479 -1828
rect 1513 -1862 1547 -1828
rect 1581 -1862 1615 -1828
rect 1649 -1862 1683 -1828
rect 1717 -1862 1751 -1828
rect 1785 -1862 1819 -1828
rect 1853 -1862 1887 -1828
rect 1921 -1862 1955 -1828
rect 1989 -1862 2023 -1828
rect 2057 -1862 2091 -1828
rect 2125 -1862 2159 -1828
rect 2193 -1862 2227 -1828
rect 2261 -1862 2295 -1828
rect 2329 -1862 2363 -1828
rect 2397 -1862 2431 -1828
rect 2465 -1862 2499 -1828
rect 2533 -1862 2567 -1828
rect 2601 -1862 2635 -1828
rect 2669 -1862 2703 -1828
rect 2737 -1862 2771 -1828
rect 2805 -1862 2839 -1828
rect 2873 -1862 2907 -1828
rect 2941 -1862 2975 -1828
rect 3009 -1862 3043 -1828
rect 3077 -1862 3111 -1828
rect 3145 -1862 3179 -1828
rect 3213 -1862 3247 -1828
rect 3281 -1862 3315 -1828
rect 3349 -1862 3383 -1828
rect 3417 -1862 3451 -1828
rect 3485 -1862 3519 -1828
rect 3553 -1862 3587 -1828
rect 3621 -1862 3655 -1828
rect 3689 -1862 3723 -1828
rect 3757 -1862 3791 -1828
rect 3825 -1862 3859 -1828
rect 3893 -1862 3927 -1828
rect 3961 -1862 4059 -1828
<< viali >>
rect -3913 1318 -3807 1712
rect -3527 1318 -3421 1712
rect -3141 1318 -3035 1712
rect -2755 1318 -2649 1712
rect -2369 1318 -2263 1712
rect -1983 1318 -1877 1712
rect -1597 1318 -1491 1712
rect -1211 1318 -1105 1712
rect -825 1318 -719 1712
rect -439 1318 -333 1712
rect -53 1318 53 1712
rect 333 1318 439 1712
rect 719 1318 825 1712
rect 1105 1318 1211 1712
rect 1491 1318 1597 1712
rect 1877 1318 1983 1712
rect 2263 1318 2369 1712
rect 2649 1318 2755 1712
rect 3035 1318 3141 1712
rect 3421 1318 3527 1712
rect 3807 1318 3913 1712
rect -3913 -1713 -3807 -1319
rect -3527 -1713 -3421 -1319
rect -3141 -1713 -3035 -1319
rect -2755 -1713 -2649 -1319
rect -2369 -1713 -2263 -1319
rect -1983 -1713 -1877 -1319
rect -1597 -1713 -1491 -1319
rect -1211 -1713 -1105 -1319
rect -825 -1713 -719 -1319
rect -439 -1713 -333 -1319
rect -53 -1713 53 -1319
rect 333 -1713 439 -1319
rect 719 -1713 825 -1319
rect 1105 -1713 1211 -1319
rect 1491 -1713 1597 -1319
rect 1877 -1713 1983 -1319
rect 2263 -1713 2369 -1319
rect 2649 -1713 2755 -1319
rect 3035 -1713 3141 -1319
rect 3421 -1713 3527 -1319
rect 3807 -1713 3913 -1319
<< metal1 >>
rect -3919 1712 -3801 1726
rect -3919 1318 -3913 1712
rect -3807 1318 -3801 1712
rect -3919 1305 -3801 1318
rect -3533 1712 -3415 1726
rect -3533 1318 -3527 1712
rect -3421 1318 -3415 1712
rect -3533 1305 -3415 1318
rect -3147 1712 -3029 1726
rect -3147 1318 -3141 1712
rect -3035 1318 -3029 1712
rect -3147 1305 -3029 1318
rect -2761 1712 -2643 1726
rect -2761 1318 -2755 1712
rect -2649 1318 -2643 1712
rect -2761 1305 -2643 1318
rect -2375 1712 -2257 1726
rect -2375 1318 -2369 1712
rect -2263 1318 -2257 1712
rect -2375 1305 -2257 1318
rect -1989 1712 -1871 1726
rect -1989 1318 -1983 1712
rect -1877 1318 -1871 1712
rect -1989 1305 -1871 1318
rect -1603 1712 -1485 1726
rect -1603 1318 -1597 1712
rect -1491 1318 -1485 1712
rect -1603 1305 -1485 1318
rect -1217 1712 -1099 1726
rect -1217 1318 -1211 1712
rect -1105 1318 -1099 1712
rect -1217 1305 -1099 1318
rect -831 1712 -713 1726
rect -831 1318 -825 1712
rect -719 1318 -713 1712
rect -831 1305 -713 1318
rect -445 1712 -327 1726
rect -445 1318 -439 1712
rect -333 1318 -327 1712
rect -445 1305 -327 1318
rect -59 1712 59 1726
rect -59 1318 -53 1712
rect 53 1318 59 1712
rect -59 1305 59 1318
rect 327 1712 445 1726
rect 327 1318 333 1712
rect 439 1318 445 1712
rect 327 1305 445 1318
rect 713 1712 831 1726
rect 713 1318 719 1712
rect 825 1318 831 1712
rect 713 1305 831 1318
rect 1099 1712 1217 1726
rect 1099 1318 1105 1712
rect 1211 1318 1217 1712
rect 1099 1305 1217 1318
rect 1485 1712 1603 1726
rect 1485 1318 1491 1712
rect 1597 1318 1603 1712
rect 1485 1305 1603 1318
rect 1871 1712 1989 1726
rect 1871 1318 1877 1712
rect 1983 1318 1989 1712
rect 1871 1305 1989 1318
rect 2257 1712 2375 1726
rect 2257 1318 2263 1712
rect 2369 1318 2375 1712
rect 2257 1305 2375 1318
rect 2643 1712 2761 1726
rect 2643 1318 2649 1712
rect 2755 1318 2761 1712
rect 2643 1305 2761 1318
rect 3029 1712 3147 1726
rect 3029 1318 3035 1712
rect 3141 1318 3147 1712
rect 3029 1305 3147 1318
rect 3415 1712 3533 1726
rect 3415 1318 3421 1712
rect 3527 1318 3533 1712
rect 3415 1305 3533 1318
rect 3801 1712 3919 1726
rect 3801 1318 3807 1712
rect 3913 1318 3919 1712
rect 3801 1305 3919 1318
rect -3919 -1319 -3801 -1305
rect -3919 -1713 -3913 -1319
rect -3807 -1713 -3801 -1319
rect -3919 -1726 -3801 -1713
rect -3533 -1319 -3415 -1305
rect -3533 -1713 -3527 -1319
rect -3421 -1713 -3415 -1319
rect -3533 -1726 -3415 -1713
rect -3147 -1319 -3029 -1305
rect -3147 -1713 -3141 -1319
rect -3035 -1713 -3029 -1319
rect -3147 -1726 -3029 -1713
rect -2761 -1319 -2643 -1305
rect -2761 -1713 -2755 -1319
rect -2649 -1713 -2643 -1319
rect -2761 -1726 -2643 -1713
rect -2375 -1319 -2257 -1305
rect -2375 -1713 -2369 -1319
rect -2263 -1713 -2257 -1319
rect -2375 -1726 -2257 -1713
rect -1989 -1319 -1871 -1305
rect -1989 -1713 -1983 -1319
rect -1877 -1713 -1871 -1319
rect -1989 -1726 -1871 -1713
rect -1603 -1319 -1485 -1305
rect -1603 -1713 -1597 -1319
rect -1491 -1713 -1485 -1319
rect -1603 -1726 -1485 -1713
rect -1217 -1319 -1099 -1305
rect -1217 -1713 -1211 -1319
rect -1105 -1713 -1099 -1319
rect -1217 -1726 -1099 -1713
rect -831 -1319 -713 -1305
rect -831 -1713 -825 -1319
rect -719 -1713 -713 -1319
rect -831 -1726 -713 -1713
rect -445 -1319 -327 -1305
rect -445 -1713 -439 -1319
rect -333 -1713 -327 -1319
rect -445 -1726 -327 -1713
rect -59 -1319 59 -1305
rect -59 -1713 -53 -1319
rect 53 -1713 59 -1319
rect -59 -1726 59 -1713
rect 327 -1319 445 -1305
rect 327 -1713 333 -1319
rect 439 -1713 445 -1319
rect 327 -1726 445 -1713
rect 713 -1319 831 -1305
rect 713 -1713 719 -1319
rect 825 -1713 831 -1319
rect 713 -1726 831 -1713
rect 1099 -1319 1217 -1305
rect 1099 -1713 1105 -1319
rect 1211 -1713 1217 -1319
rect 1099 -1726 1217 -1713
rect 1485 -1319 1603 -1305
rect 1485 -1713 1491 -1319
rect 1597 -1713 1603 -1319
rect 1485 -1726 1603 -1713
rect 1871 -1319 1989 -1305
rect 1871 -1713 1877 -1319
rect 1983 -1713 1989 -1319
rect 1871 -1726 1989 -1713
rect 2257 -1319 2375 -1305
rect 2257 -1713 2263 -1319
rect 2369 -1713 2375 -1319
rect 2257 -1726 2375 -1713
rect 2643 -1319 2761 -1305
rect 2643 -1713 2649 -1319
rect 2755 -1713 2761 -1319
rect 2643 -1726 2761 -1713
rect 3029 -1319 3147 -1305
rect 3029 -1713 3035 -1319
rect 3141 -1713 3147 -1319
rect 3029 -1726 3147 -1713
rect 3415 -1319 3533 -1305
rect 3415 -1713 3421 -1319
rect 3527 -1713 3533 -1319
rect 3415 -1726 3533 -1713
rect 3801 -1319 3919 -1305
rect 3801 -1713 3807 -1319
rect 3913 -1713 3919 -1319
rect 3801 -1726 3919 -1713
<< properties >>
string FIXED_BBOX -4042 -1845 4042 1845
<< end >>
