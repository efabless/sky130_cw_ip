magic
tech sky130A
magscale 1 2
timestamp 1715625863
<< pwell >>
rect -26184 8606 -13334 8692
rect -26184 5351 -26098 8606
rect -13420 5351 -13334 8606
rect -26184 5265 -13334 5351
<< psubdiff >>
rect -26158 8632 -26000 8666
rect -25966 8632 -25932 8666
rect -25898 8632 -25864 8666
rect -25830 8632 -25796 8666
rect -25762 8632 -25728 8666
rect -25694 8632 -25660 8666
rect -25626 8632 -25592 8666
rect -25558 8632 -25524 8666
rect -25490 8632 -25456 8666
rect -25422 8632 -25388 8666
rect -25354 8632 -25320 8666
rect -25286 8632 -25252 8666
rect -25218 8632 -25184 8666
rect -25150 8632 -25116 8666
rect -25082 8632 -25048 8666
rect -25014 8632 -24980 8666
rect -24946 8632 -24912 8666
rect -24878 8632 -24844 8666
rect -24810 8632 -24776 8666
rect -24742 8632 -24708 8666
rect -24674 8632 -24640 8666
rect -24606 8632 -24572 8666
rect -24538 8632 -24504 8666
rect -24470 8632 -24436 8666
rect -24402 8632 -24368 8666
rect -24334 8632 -24300 8666
rect -24266 8632 -24232 8666
rect -24198 8632 -24164 8666
rect -24130 8632 -24096 8666
rect -24062 8632 -24028 8666
rect -23994 8632 -23960 8666
rect -23926 8632 -23892 8666
rect -23858 8632 -23824 8666
rect -23790 8632 -23756 8666
rect -23722 8632 -23688 8666
rect -23654 8632 -23620 8666
rect -23586 8632 -23552 8666
rect -23518 8632 -23484 8666
rect -23450 8632 -23416 8666
rect -23382 8632 -23348 8666
rect -23314 8632 -23280 8666
rect -23246 8632 -23212 8666
rect -23178 8632 -23144 8666
rect -23110 8632 -23076 8666
rect -23042 8632 -23008 8666
rect -22974 8632 -22940 8666
rect -22906 8632 -22872 8666
rect -22838 8632 -22804 8666
rect -22770 8632 -22736 8666
rect -22702 8632 -22668 8666
rect -22634 8632 -22600 8666
rect -22566 8632 -22532 8666
rect -22498 8632 -22464 8666
rect -22430 8632 -22396 8666
rect -22362 8632 -22328 8666
rect -22294 8632 -22260 8666
rect -22226 8632 -22192 8666
rect -22158 8632 -22124 8666
rect -22090 8632 -22056 8666
rect -22022 8632 -21988 8666
rect -21954 8632 -21920 8666
rect -21886 8632 -21852 8666
rect -21818 8632 -21784 8666
rect -21750 8632 -21716 8666
rect -21682 8632 -21648 8666
rect -21614 8632 -21580 8666
rect -21546 8632 -21512 8666
rect -21478 8632 -21444 8666
rect -21410 8632 -21376 8666
rect -21342 8632 -21308 8666
rect -21274 8632 -21240 8666
rect -21206 8632 -21172 8666
rect -21138 8632 -21104 8666
rect -21070 8632 -21036 8666
rect -21002 8632 -20968 8666
rect -20934 8632 -20900 8666
rect -20866 8632 -20832 8666
rect -20798 8632 -20764 8666
rect -20730 8632 -20696 8666
rect -20662 8632 -20628 8666
rect -20594 8632 -20560 8666
rect -20526 8632 -20492 8666
rect -20458 8632 -20424 8666
rect -20390 8632 -20356 8666
rect -20322 8632 -20288 8666
rect -20254 8632 -20220 8666
rect -20186 8632 -20152 8666
rect -20118 8632 -20084 8666
rect -20050 8632 -20016 8666
rect -19982 8632 -19948 8666
rect -19914 8632 -19880 8666
rect -19846 8632 -19812 8666
rect -19778 8632 -19744 8666
rect -19710 8632 -19676 8666
rect -19642 8632 -19608 8666
rect -19574 8632 -19540 8666
rect -19506 8632 -19472 8666
rect -19438 8632 -19404 8666
rect -19370 8632 -19336 8666
rect -19302 8632 -19268 8666
rect -19234 8632 -19200 8666
rect -19166 8632 -19132 8666
rect -19098 8632 -19064 8666
rect -19030 8632 -18996 8666
rect -18962 8632 -18928 8666
rect -18894 8632 -18860 8666
rect -18826 8632 -18792 8666
rect -18758 8632 -18724 8666
rect -18690 8632 -18656 8666
rect -18622 8632 -18588 8666
rect -18554 8632 -18520 8666
rect -18486 8632 -18452 8666
rect -18418 8632 -18384 8666
rect -18350 8632 -18316 8666
rect -18282 8632 -18248 8666
rect -18214 8632 -18180 8666
rect -18146 8632 -18112 8666
rect -18078 8632 -18044 8666
rect -18010 8632 -17976 8666
rect -17942 8632 -17908 8666
rect -17874 8632 -17840 8666
rect -17806 8632 -17772 8666
rect -17738 8632 -17704 8666
rect -17670 8632 -17636 8666
rect -17602 8632 -17568 8666
rect -17534 8632 -17500 8666
rect -17466 8632 -17432 8666
rect -17398 8632 -17364 8666
rect -17330 8632 -17296 8666
rect -17262 8632 -17228 8666
rect -17194 8632 -17160 8666
rect -17126 8632 -17092 8666
rect -17058 8632 -17024 8666
rect -16990 8632 -16956 8666
rect -16922 8632 -16888 8666
rect -16854 8632 -16820 8666
rect -16786 8632 -16752 8666
rect -16718 8632 -16684 8666
rect -16650 8632 -16616 8666
rect -16582 8632 -16548 8666
rect -16514 8632 -16480 8666
rect -16446 8632 -16412 8666
rect -16378 8632 -16344 8666
rect -16310 8632 -16276 8666
rect -16242 8632 -16208 8666
rect -16174 8632 -16140 8666
rect -16106 8632 -16072 8666
rect -16038 8632 -16004 8666
rect -15970 8632 -15936 8666
rect -15902 8632 -15868 8666
rect -15834 8632 -15800 8666
rect -15766 8632 -15732 8666
rect -15698 8632 -15664 8666
rect -15630 8632 -15596 8666
rect -15562 8632 -15528 8666
rect -15494 8632 -15460 8666
rect -15426 8632 -15392 8666
rect -15358 8632 -15324 8666
rect -15290 8632 -15256 8666
rect -15222 8632 -15188 8666
rect -15154 8632 -15120 8666
rect -15086 8632 -15052 8666
rect -15018 8632 -14984 8666
rect -14950 8632 -14916 8666
rect -14882 8632 -14848 8666
rect -14814 8632 -14780 8666
rect -14746 8632 -14712 8666
rect -14678 8632 -14644 8666
rect -14610 8632 -14576 8666
rect -14542 8632 -14508 8666
rect -14474 8632 -14440 8666
rect -14406 8632 -14372 8666
rect -14338 8632 -14304 8666
rect -14270 8632 -14236 8666
rect -14202 8632 -14168 8666
rect -14134 8632 -14100 8666
rect -14066 8632 -14032 8666
rect -13998 8632 -13964 8666
rect -13930 8632 -13896 8666
rect -13862 8632 -13828 8666
rect -13794 8632 -13760 8666
rect -13726 8632 -13692 8666
rect -13658 8632 -13624 8666
rect -13590 8632 -13360 8666
rect -26158 8466 -26124 8632
rect -26158 8398 -26124 8432
rect -26158 8330 -26124 8364
rect -26158 8262 -26124 8296
rect -26158 8194 -26124 8228
rect -26158 8126 -26124 8160
rect -26158 8058 -26124 8092
rect -26158 7990 -26124 8024
rect -26158 7922 -26124 7956
rect -26158 7854 -26124 7888
rect -26158 7786 -26124 7820
rect -26158 7718 -26124 7752
rect -26158 7650 -26124 7684
rect -26158 7582 -26124 7616
rect -26158 7514 -26124 7548
rect -26158 7446 -26124 7480
rect -26158 7378 -26124 7412
rect -26158 7310 -26124 7344
rect -26158 7242 -26124 7276
rect -26158 7174 -26124 7208
rect -26158 7106 -26124 7140
rect -26158 7038 -26124 7072
rect -26158 6970 -26124 7004
rect -26158 6902 -26124 6936
rect -26158 6834 -26124 6868
rect -26158 6766 -26124 6800
rect -26158 6698 -26124 6732
rect -26158 6630 -26124 6664
rect -26158 6562 -26124 6596
rect -26158 6494 -26124 6528
rect -26158 6426 -26124 6460
rect -26158 6358 -26124 6392
rect -26158 6290 -26124 6324
rect -26158 6222 -26124 6256
rect -26158 6154 -26124 6188
rect -26158 6086 -26124 6120
rect -26158 6018 -26124 6052
rect -26158 5950 -26124 5984
rect -26158 5882 -26124 5916
rect -26158 5814 -26124 5848
rect -26158 5746 -26124 5780
rect -26158 5678 -26124 5712
rect -26158 5610 -26124 5644
rect -26158 5542 -26124 5576
rect -26158 5325 -26124 5508
rect -13394 8466 -13360 8632
rect -13394 8398 -13360 8432
rect -13394 8330 -13360 8364
rect -13394 8262 -13360 8296
rect -13394 8194 -13360 8228
rect -13394 8126 -13360 8160
rect -13394 8058 -13360 8092
rect -13394 7990 -13360 8024
rect -13394 7922 -13360 7956
rect -13394 7854 -13360 7888
rect -13394 7786 -13360 7820
rect -13394 7718 -13360 7752
rect -13394 7650 -13360 7684
rect -13394 7582 -13360 7616
rect -13394 7514 -13360 7548
rect -13394 7446 -13360 7480
rect -13394 7378 -13360 7412
rect -13394 7310 -13360 7344
rect -13394 7242 -13360 7276
rect -13394 7174 -13360 7208
rect -13394 7106 -13360 7140
rect -13394 7038 -13360 7072
rect -13394 6970 -13360 7004
rect -13394 6902 -13360 6936
rect -13394 6834 -13360 6868
rect -13394 6766 -13360 6800
rect -13394 6698 -13360 6732
rect -13394 6630 -13360 6664
rect -13394 6562 -13360 6596
rect -13394 6494 -13360 6528
rect -13394 6426 -13360 6460
rect -13394 6358 -13360 6392
rect -13394 6290 -13360 6324
rect -13394 6222 -13360 6256
rect -13394 6154 -13360 6188
rect -13394 6086 -13360 6120
rect -13394 6018 -13360 6052
rect -13394 5950 -13360 5984
rect -13394 5882 -13360 5916
rect -13394 5814 -13360 5848
rect -13394 5746 -13360 5780
rect -13394 5678 -13360 5712
rect -13394 5610 -13360 5644
rect -13394 5542 -13360 5576
rect -13394 5325 -13360 5508
rect -26158 5291 -25958 5325
rect -25924 5291 -25890 5325
rect -25856 5291 -25822 5325
rect -25788 5291 -25754 5325
rect -25720 5291 -25686 5325
rect -25652 5291 -25618 5325
rect -25584 5291 -25550 5325
rect -25516 5291 -25482 5325
rect -25448 5291 -25414 5325
rect -25380 5291 -25346 5325
rect -25312 5291 -25278 5325
rect -25244 5291 -25210 5325
rect -25176 5291 -25142 5325
rect -25108 5291 -25074 5325
rect -25040 5291 -25006 5325
rect -24972 5291 -24938 5325
rect -24904 5291 -24870 5325
rect -24836 5291 -24802 5325
rect -24768 5291 -24734 5325
rect -24700 5291 -24666 5325
rect -24632 5291 -24598 5325
rect -24564 5291 -24530 5325
rect -24496 5291 -24462 5325
rect -24428 5291 -24394 5325
rect -24360 5291 -24326 5325
rect -24292 5291 -24258 5325
rect -24224 5291 -24190 5325
rect -24156 5291 -24122 5325
rect -24088 5291 -24054 5325
rect -24020 5291 -23986 5325
rect -23952 5291 -23918 5325
rect -23884 5291 -23850 5325
rect -23816 5291 -23782 5325
rect -23748 5291 -23714 5325
rect -23680 5291 -23646 5325
rect -23612 5291 -23578 5325
rect -23544 5291 -23510 5325
rect -23476 5291 -23442 5325
rect -23408 5291 -23374 5325
rect -23340 5291 -23306 5325
rect -23272 5291 -23238 5325
rect -23204 5291 -23170 5325
rect -23136 5291 -23102 5325
rect -23068 5291 -23034 5325
rect -23000 5291 -22966 5325
rect -22932 5291 -22898 5325
rect -22864 5291 -22830 5325
rect -22796 5291 -22762 5325
rect -22728 5291 -22694 5325
rect -22660 5291 -22626 5325
rect -22592 5291 -22558 5325
rect -22524 5291 -22490 5325
rect -22456 5291 -22422 5325
rect -22388 5291 -22354 5325
rect -22320 5291 -22286 5325
rect -22252 5291 -22218 5325
rect -22184 5291 -22150 5325
rect -22116 5291 -22082 5325
rect -22048 5291 -22014 5325
rect -21980 5291 -21946 5325
rect -21912 5291 -21878 5325
rect -21844 5291 -21810 5325
rect -21776 5291 -21742 5325
rect -21708 5291 -21674 5325
rect -21640 5291 -21606 5325
rect -21572 5291 -21538 5325
rect -21504 5291 -21470 5325
rect -21436 5291 -21402 5325
rect -21368 5291 -21334 5325
rect -21300 5291 -21266 5325
rect -21232 5291 -21198 5325
rect -21164 5291 -21130 5325
rect -21096 5291 -21062 5325
rect -21028 5291 -20994 5325
rect -20960 5291 -20926 5325
rect -20892 5291 -20858 5325
rect -20824 5291 -20790 5325
rect -20756 5291 -20722 5325
rect -20688 5291 -20654 5325
rect -20620 5291 -20586 5325
rect -20552 5291 -20518 5325
rect -20484 5291 -20450 5325
rect -20416 5291 -20382 5325
rect -20348 5291 -20314 5325
rect -20280 5291 -20246 5325
rect -20212 5291 -20178 5325
rect -20144 5291 -20110 5325
rect -20076 5291 -20042 5325
rect -20008 5291 -19974 5325
rect -19940 5291 -19906 5325
rect -19872 5291 -19838 5325
rect -19804 5291 -19770 5325
rect -19736 5291 -19702 5325
rect -19668 5291 -19634 5325
rect -19600 5291 -19566 5325
rect -19532 5291 -19498 5325
rect -19464 5291 -19430 5325
rect -19396 5291 -19362 5325
rect -19328 5291 -19294 5325
rect -19260 5291 -19226 5325
rect -19192 5291 -19158 5325
rect -19124 5291 -19090 5325
rect -19056 5291 -19022 5325
rect -18988 5291 -18954 5325
rect -18920 5291 -18886 5325
rect -18852 5291 -18818 5325
rect -18784 5291 -18750 5325
rect -18716 5291 -18682 5325
rect -18648 5291 -18614 5325
rect -18580 5291 -18546 5325
rect -18512 5291 -18478 5325
rect -18444 5291 -18410 5325
rect -18376 5291 -18342 5325
rect -18308 5291 -18274 5325
rect -18240 5291 -18206 5325
rect -18172 5291 -18138 5325
rect -18104 5291 -18070 5325
rect -18036 5291 -18002 5325
rect -17968 5291 -17934 5325
rect -17900 5291 -17866 5325
rect -17832 5291 -17798 5325
rect -17764 5291 -17730 5325
rect -17696 5291 -17662 5325
rect -17628 5291 -17594 5325
rect -17560 5291 -17526 5325
rect -17492 5291 -17458 5325
rect -17424 5291 -17390 5325
rect -17356 5291 -17322 5325
rect -17288 5291 -17254 5325
rect -17220 5291 -17186 5325
rect -17152 5291 -17118 5325
rect -17084 5291 -17050 5325
rect -17016 5291 -16982 5325
rect -16948 5291 -16914 5325
rect -16880 5291 -16846 5325
rect -16812 5291 -16778 5325
rect -16744 5291 -16710 5325
rect -16676 5291 -16642 5325
rect -16608 5291 -16574 5325
rect -16540 5291 -16506 5325
rect -16472 5291 -16438 5325
rect -16404 5291 -16370 5325
rect -16336 5291 -16302 5325
rect -16268 5291 -16234 5325
rect -16200 5291 -16166 5325
rect -16132 5291 -16098 5325
rect -16064 5291 -16030 5325
rect -15996 5291 -15962 5325
rect -15928 5291 -15894 5325
rect -15860 5291 -15826 5325
rect -15792 5291 -15758 5325
rect -15724 5291 -15690 5325
rect -15656 5291 -15622 5325
rect -15588 5291 -15554 5325
rect -15520 5291 -15486 5325
rect -15452 5291 -15418 5325
rect -15384 5291 -15350 5325
rect -15316 5291 -15282 5325
rect -15248 5291 -15214 5325
rect -15180 5291 -15146 5325
rect -15112 5291 -15078 5325
rect -15044 5291 -15010 5325
rect -14976 5291 -14942 5325
rect -14908 5291 -14874 5325
rect -14840 5291 -14806 5325
rect -14772 5291 -14738 5325
rect -14704 5291 -14670 5325
rect -14636 5291 -14602 5325
rect -14568 5291 -14534 5325
rect -14500 5291 -14466 5325
rect -14432 5291 -14398 5325
rect -14364 5291 -14330 5325
rect -14296 5291 -14262 5325
rect -14228 5291 -14194 5325
rect -14160 5291 -14126 5325
rect -14092 5291 -14058 5325
rect -14024 5291 -13990 5325
rect -13956 5291 -13922 5325
rect -13888 5291 -13854 5325
rect -13820 5291 -13786 5325
rect -13752 5291 -13718 5325
rect -13684 5291 -13650 5325
rect -13616 5291 -13360 5325
<< psubdiffcont >>
rect -26000 8632 -25966 8666
rect -25932 8632 -25898 8666
rect -25864 8632 -25830 8666
rect -25796 8632 -25762 8666
rect -25728 8632 -25694 8666
rect -25660 8632 -25626 8666
rect -25592 8632 -25558 8666
rect -25524 8632 -25490 8666
rect -25456 8632 -25422 8666
rect -25388 8632 -25354 8666
rect -25320 8632 -25286 8666
rect -25252 8632 -25218 8666
rect -25184 8632 -25150 8666
rect -25116 8632 -25082 8666
rect -25048 8632 -25014 8666
rect -24980 8632 -24946 8666
rect -24912 8632 -24878 8666
rect -24844 8632 -24810 8666
rect -24776 8632 -24742 8666
rect -24708 8632 -24674 8666
rect -24640 8632 -24606 8666
rect -24572 8632 -24538 8666
rect -24504 8632 -24470 8666
rect -24436 8632 -24402 8666
rect -24368 8632 -24334 8666
rect -24300 8632 -24266 8666
rect -24232 8632 -24198 8666
rect -24164 8632 -24130 8666
rect -24096 8632 -24062 8666
rect -24028 8632 -23994 8666
rect -23960 8632 -23926 8666
rect -23892 8632 -23858 8666
rect -23824 8632 -23790 8666
rect -23756 8632 -23722 8666
rect -23688 8632 -23654 8666
rect -23620 8632 -23586 8666
rect -23552 8632 -23518 8666
rect -23484 8632 -23450 8666
rect -23416 8632 -23382 8666
rect -23348 8632 -23314 8666
rect -23280 8632 -23246 8666
rect -23212 8632 -23178 8666
rect -23144 8632 -23110 8666
rect -23076 8632 -23042 8666
rect -23008 8632 -22974 8666
rect -22940 8632 -22906 8666
rect -22872 8632 -22838 8666
rect -22804 8632 -22770 8666
rect -22736 8632 -22702 8666
rect -22668 8632 -22634 8666
rect -22600 8632 -22566 8666
rect -22532 8632 -22498 8666
rect -22464 8632 -22430 8666
rect -22396 8632 -22362 8666
rect -22328 8632 -22294 8666
rect -22260 8632 -22226 8666
rect -22192 8632 -22158 8666
rect -22124 8632 -22090 8666
rect -22056 8632 -22022 8666
rect -21988 8632 -21954 8666
rect -21920 8632 -21886 8666
rect -21852 8632 -21818 8666
rect -21784 8632 -21750 8666
rect -21716 8632 -21682 8666
rect -21648 8632 -21614 8666
rect -21580 8632 -21546 8666
rect -21512 8632 -21478 8666
rect -21444 8632 -21410 8666
rect -21376 8632 -21342 8666
rect -21308 8632 -21274 8666
rect -21240 8632 -21206 8666
rect -21172 8632 -21138 8666
rect -21104 8632 -21070 8666
rect -21036 8632 -21002 8666
rect -20968 8632 -20934 8666
rect -20900 8632 -20866 8666
rect -20832 8632 -20798 8666
rect -20764 8632 -20730 8666
rect -20696 8632 -20662 8666
rect -20628 8632 -20594 8666
rect -20560 8632 -20526 8666
rect -20492 8632 -20458 8666
rect -20424 8632 -20390 8666
rect -20356 8632 -20322 8666
rect -20288 8632 -20254 8666
rect -20220 8632 -20186 8666
rect -20152 8632 -20118 8666
rect -20084 8632 -20050 8666
rect -20016 8632 -19982 8666
rect -19948 8632 -19914 8666
rect -19880 8632 -19846 8666
rect -19812 8632 -19778 8666
rect -19744 8632 -19710 8666
rect -19676 8632 -19642 8666
rect -19608 8632 -19574 8666
rect -19540 8632 -19506 8666
rect -19472 8632 -19438 8666
rect -19404 8632 -19370 8666
rect -19336 8632 -19302 8666
rect -19268 8632 -19234 8666
rect -19200 8632 -19166 8666
rect -19132 8632 -19098 8666
rect -19064 8632 -19030 8666
rect -18996 8632 -18962 8666
rect -18928 8632 -18894 8666
rect -18860 8632 -18826 8666
rect -18792 8632 -18758 8666
rect -18724 8632 -18690 8666
rect -18656 8632 -18622 8666
rect -18588 8632 -18554 8666
rect -18520 8632 -18486 8666
rect -18452 8632 -18418 8666
rect -18384 8632 -18350 8666
rect -18316 8632 -18282 8666
rect -18248 8632 -18214 8666
rect -18180 8632 -18146 8666
rect -18112 8632 -18078 8666
rect -18044 8632 -18010 8666
rect -17976 8632 -17942 8666
rect -17908 8632 -17874 8666
rect -17840 8632 -17806 8666
rect -17772 8632 -17738 8666
rect -17704 8632 -17670 8666
rect -17636 8632 -17602 8666
rect -17568 8632 -17534 8666
rect -17500 8632 -17466 8666
rect -17432 8632 -17398 8666
rect -17364 8632 -17330 8666
rect -17296 8632 -17262 8666
rect -17228 8632 -17194 8666
rect -17160 8632 -17126 8666
rect -17092 8632 -17058 8666
rect -17024 8632 -16990 8666
rect -16956 8632 -16922 8666
rect -16888 8632 -16854 8666
rect -16820 8632 -16786 8666
rect -16752 8632 -16718 8666
rect -16684 8632 -16650 8666
rect -16616 8632 -16582 8666
rect -16548 8632 -16514 8666
rect -16480 8632 -16446 8666
rect -16412 8632 -16378 8666
rect -16344 8632 -16310 8666
rect -16276 8632 -16242 8666
rect -16208 8632 -16174 8666
rect -16140 8632 -16106 8666
rect -16072 8632 -16038 8666
rect -16004 8632 -15970 8666
rect -15936 8632 -15902 8666
rect -15868 8632 -15834 8666
rect -15800 8632 -15766 8666
rect -15732 8632 -15698 8666
rect -15664 8632 -15630 8666
rect -15596 8632 -15562 8666
rect -15528 8632 -15494 8666
rect -15460 8632 -15426 8666
rect -15392 8632 -15358 8666
rect -15324 8632 -15290 8666
rect -15256 8632 -15222 8666
rect -15188 8632 -15154 8666
rect -15120 8632 -15086 8666
rect -15052 8632 -15018 8666
rect -14984 8632 -14950 8666
rect -14916 8632 -14882 8666
rect -14848 8632 -14814 8666
rect -14780 8632 -14746 8666
rect -14712 8632 -14678 8666
rect -14644 8632 -14610 8666
rect -14576 8632 -14542 8666
rect -14508 8632 -14474 8666
rect -14440 8632 -14406 8666
rect -14372 8632 -14338 8666
rect -14304 8632 -14270 8666
rect -14236 8632 -14202 8666
rect -14168 8632 -14134 8666
rect -14100 8632 -14066 8666
rect -14032 8632 -13998 8666
rect -13964 8632 -13930 8666
rect -13896 8632 -13862 8666
rect -13828 8632 -13794 8666
rect -13760 8632 -13726 8666
rect -13692 8632 -13658 8666
rect -13624 8632 -13590 8666
rect -26158 8432 -26124 8466
rect -26158 8364 -26124 8398
rect -26158 8296 -26124 8330
rect -26158 8228 -26124 8262
rect -26158 8160 -26124 8194
rect -26158 8092 -26124 8126
rect -26158 8024 -26124 8058
rect -26158 7956 -26124 7990
rect -26158 7888 -26124 7922
rect -26158 7820 -26124 7854
rect -26158 7752 -26124 7786
rect -26158 7684 -26124 7718
rect -26158 7616 -26124 7650
rect -26158 7548 -26124 7582
rect -26158 7480 -26124 7514
rect -26158 7412 -26124 7446
rect -26158 7344 -26124 7378
rect -26158 7276 -26124 7310
rect -26158 7208 -26124 7242
rect -26158 7140 -26124 7174
rect -26158 7072 -26124 7106
rect -26158 7004 -26124 7038
rect -26158 6936 -26124 6970
rect -26158 6868 -26124 6902
rect -26158 6800 -26124 6834
rect -26158 6732 -26124 6766
rect -26158 6664 -26124 6698
rect -26158 6596 -26124 6630
rect -26158 6528 -26124 6562
rect -26158 6460 -26124 6494
rect -26158 6392 -26124 6426
rect -26158 6324 -26124 6358
rect -26158 6256 -26124 6290
rect -26158 6188 -26124 6222
rect -26158 6120 -26124 6154
rect -26158 6052 -26124 6086
rect -26158 5984 -26124 6018
rect -26158 5916 -26124 5950
rect -26158 5848 -26124 5882
rect -26158 5780 -26124 5814
rect -26158 5712 -26124 5746
rect -26158 5644 -26124 5678
rect -26158 5576 -26124 5610
rect -26158 5508 -26124 5542
rect -13394 8432 -13360 8466
rect -13394 8364 -13360 8398
rect -13394 8296 -13360 8330
rect -13394 8228 -13360 8262
rect -13394 8160 -13360 8194
rect -13394 8092 -13360 8126
rect -13394 8024 -13360 8058
rect -13394 7956 -13360 7990
rect -13394 7888 -13360 7922
rect -13394 7820 -13360 7854
rect -13394 7752 -13360 7786
rect -13394 7684 -13360 7718
rect -13394 7616 -13360 7650
rect -13394 7548 -13360 7582
rect -13394 7480 -13360 7514
rect -13394 7412 -13360 7446
rect -13394 7344 -13360 7378
rect -13394 7276 -13360 7310
rect -13394 7208 -13360 7242
rect -13394 7140 -13360 7174
rect -13394 7072 -13360 7106
rect -13394 7004 -13360 7038
rect -13394 6936 -13360 6970
rect -13394 6868 -13360 6902
rect -13394 6800 -13360 6834
rect -13394 6732 -13360 6766
rect -13394 6664 -13360 6698
rect -13394 6596 -13360 6630
rect -13394 6528 -13360 6562
rect -13394 6460 -13360 6494
rect -13394 6392 -13360 6426
rect -13394 6324 -13360 6358
rect -13394 6256 -13360 6290
rect -13394 6188 -13360 6222
rect -13394 6120 -13360 6154
rect -13394 6052 -13360 6086
rect -13394 5984 -13360 6018
rect -13394 5916 -13360 5950
rect -13394 5848 -13360 5882
rect -13394 5780 -13360 5814
rect -13394 5712 -13360 5746
rect -13394 5644 -13360 5678
rect -13394 5576 -13360 5610
rect -13394 5508 -13360 5542
rect -25958 5291 -25924 5325
rect -25890 5291 -25856 5325
rect -25822 5291 -25788 5325
rect -25754 5291 -25720 5325
rect -25686 5291 -25652 5325
rect -25618 5291 -25584 5325
rect -25550 5291 -25516 5325
rect -25482 5291 -25448 5325
rect -25414 5291 -25380 5325
rect -25346 5291 -25312 5325
rect -25278 5291 -25244 5325
rect -25210 5291 -25176 5325
rect -25142 5291 -25108 5325
rect -25074 5291 -25040 5325
rect -25006 5291 -24972 5325
rect -24938 5291 -24904 5325
rect -24870 5291 -24836 5325
rect -24802 5291 -24768 5325
rect -24734 5291 -24700 5325
rect -24666 5291 -24632 5325
rect -24598 5291 -24564 5325
rect -24530 5291 -24496 5325
rect -24462 5291 -24428 5325
rect -24394 5291 -24360 5325
rect -24326 5291 -24292 5325
rect -24258 5291 -24224 5325
rect -24190 5291 -24156 5325
rect -24122 5291 -24088 5325
rect -24054 5291 -24020 5325
rect -23986 5291 -23952 5325
rect -23918 5291 -23884 5325
rect -23850 5291 -23816 5325
rect -23782 5291 -23748 5325
rect -23714 5291 -23680 5325
rect -23646 5291 -23612 5325
rect -23578 5291 -23544 5325
rect -23510 5291 -23476 5325
rect -23442 5291 -23408 5325
rect -23374 5291 -23340 5325
rect -23306 5291 -23272 5325
rect -23238 5291 -23204 5325
rect -23170 5291 -23136 5325
rect -23102 5291 -23068 5325
rect -23034 5291 -23000 5325
rect -22966 5291 -22932 5325
rect -22898 5291 -22864 5325
rect -22830 5291 -22796 5325
rect -22762 5291 -22728 5325
rect -22694 5291 -22660 5325
rect -22626 5291 -22592 5325
rect -22558 5291 -22524 5325
rect -22490 5291 -22456 5325
rect -22422 5291 -22388 5325
rect -22354 5291 -22320 5325
rect -22286 5291 -22252 5325
rect -22218 5291 -22184 5325
rect -22150 5291 -22116 5325
rect -22082 5291 -22048 5325
rect -22014 5291 -21980 5325
rect -21946 5291 -21912 5325
rect -21878 5291 -21844 5325
rect -21810 5291 -21776 5325
rect -21742 5291 -21708 5325
rect -21674 5291 -21640 5325
rect -21606 5291 -21572 5325
rect -21538 5291 -21504 5325
rect -21470 5291 -21436 5325
rect -21402 5291 -21368 5325
rect -21334 5291 -21300 5325
rect -21266 5291 -21232 5325
rect -21198 5291 -21164 5325
rect -21130 5291 -21096 5325
rect -21062 5291 -21028 5325
rect -20994 5291 -20960 5325
rect -20926 5291 -20892 5325
rect -20858 5291 -20824 5325
rect -20790 5291 -20756 5325
rect -20722 5291 -20688 5325
rect -20654 5291 -20620 5325
rect -20586 5291 -20552 5325
rect -20518 5291 -20484 5325
rect -20450 5291 -20416 5325
rect -20382 5291 -20348 5325
rect -20314 5291 -20280 5325
rect -20246 5291 -20212 5325
rect -20178 5291 -20144 5325
rect -20110 5291 -20076 5325
rect -20042 5291 -20008 5325
rect -19974 5291 -19940 5325
rect -19906 5291 -19872 5325
rect -19838 5291 -19804 5325
rect -19770 5291 -19736 5325
rect -19702 5291 -19668 5325
rect -19634 5291 -19600 5325
rect -19566 5291 -19532 5325
rect -19498 5291 -19464 5325
rect -19430 5291 -19396 5325
rect -19362 5291 -19328 5325
rect -19294 5291 -19260 5325
rect -19226 5291 -19192 5325
rect -19158 5291 -19124 5325
rect -19090 5291 -19056 5325
rect -19022 5291 -18988 5325
rect -18954 5291 -18920 5325
rect -18886 5291 -18852 5325
rect -18818 5291 -18784 5325
rect -18750 5291 -18716 5325
rect -18682 5291 -18648 5325
rect -18614 5291 -18580 5325
rect -18546 5291 -18512 5325
rect -18478 5291 -18444 5325
rect -18410 5291 -18376 5325
rect -18342 5291 -18308 5325
rect -18274 5291 -18240 5325
rect -18206 5291 -18172 5325
rect -18138 5291 -18104 5325
rect -18070 5291 -18036 5325
rect -18002 5291 -17968 5325
rect -17934 5291 -17900 5325
rect -17866 5291 -17832 5325
rect -17798 5291 -17764 5325
rect -17730 5291 -17696 5325
rect -17662 5291 -17628 5325
rect -17594 5291 -17560 5325
rect -17526 5291 -17492 5325
rect -17458 5291 -17424 5325
rect -17390 5291 -17356 5325
rect -17322 5291 -17288 5325
rect -17254 5291 -17220 5325
rect -17186 5291 -17152 5325
rect -17118 5291 -17084 5325
rect -17050 5291 -17016 5325
rect -16982 5291 -16948 5325
rect -16914 5291 -16880 5325
rect -16846 5291 -16812 5325
rect -16778 5291 -16744 5325
rect -16710 5291 -16676 5325
rect -16642 5291 -16608 5325
rect -16574 5291 -16540 5325
rect -16506 5291 -16472 5325
rect -16438 5291 -16404 5325
rect -16370 5291 -16336 5325
rect -16302 5291 -16268 5325
rect -16234 5291 -16200 5325
rect -16166 5291 -16132 5325
rect -16098 5291 -16064 5325
rect -16030 5291 -15996 5325
rect -15962 5291 -15928 5325
rect -15894 5291 -15860 5325
rect -15826 5291 -15792 5325
rect -15758 5291 -15724 5325
rect -15690 5291 -15656 5325
rect -15622 5291 -15588 5325
rect -15554 5291 -15520 5325
rect -15486 5291 -15452 5325
rect -15418 5291 -15384 5325
rect -15350 5291 -15316 5325
rect -15282 5291 -15248 5325
rect -15214 5291 -15180 5325
rect -15146 5291 -15112 5325
rect -15078 5291 -15044 5325
rect -15010 5291 -14976 5325
rect -14942 5291 -14908 5325
rect -14874 5291 -14840 5325
rect -14806 5291 -14772 5325
rect -14738 5291 -14704 5325
rect -14670 5291 -14636 5325
rect -14602 5291 -14568 5325
rect -14534 5291 -14500 5325
rect -14466 5291 -14432 5325
rect -14398 5291 -14364 5325
rect -14330 5291 -14296 5325
rect -14262 5291 -14228 5325
rect -14194 5291 -14160 5325
rect -14126 5291 -14092 5325
rect -14058 5291 -14024 5325
rect -13990 5291 -13956 5325
rect -13922 5291 -13888 5325
rect -13854 5291 -13820 5325
rect -13786 5291 -13752 5325
rect -13718 5291 -13684 5325
rect -13650 5291 -13616 5325
<< locali >>
rect -26158 8632 -26000 8666
rect -25966 8632 -25932 8666
rect -25898 8632 -25864 8666
rect -25830 8632 -25796 8666
rect -25762 8632 -25728 8666
rect -25694 8632 -25660 8666
rect -25626 8632 -25592 8666
rect -25558 8632 -25524 8666
rect -25490 8632 -25456 8666
rect -25422 8632 -25388 8666
rect -25354 8632 -25320 8666
rect -25286 8632 -25252 8666
rect -25218 8632 -25184 8666
rect -25150 8632 -25116 8666
rect -25082 8632 -25048 8666
rect -25014 8632 -24980 8666
rect -24946 8632 -24912 8666
rect -24878 8632 -24844 8666
rect -24810 8632 -24776 8666
rect -24742 8632 -24708 8666
rect -24674 8632 -24640 8666
rect -24606 8632 -24572 8666
rect -24538 8632 -24504 8666
rect -24470 8632 -24436 8666
rect -24402 8632 -24368 8666
rect -24334 8632 -24300 8666
rect -24266 8632 -24232 8666
rect -24198 8632 -24164 8666
rect -24130 8632 -24096 8666
rect -24062 8632 -24028 8666
rect -23994 8632 -23960 8666
rect -23926 8632 -23892 8666
rect -23858 8632 -23824 8666
rect -23790 8632 -23756 8666
rect -23722 8632 -23688 8666
rect -23654 8632 -23620 8666
rect -23586 8632 -23552 8666
rect -23518 8632 -23484 8666
rect -23450 8632 -23416 8666
rect -23382 8632 -23348 8666
rect -23314 8632 -23280 8666
rect -23246 8632 -23212 8666
rect -23178 8632 -23144 8666
rect -23110 8632 -23076 8666
rect -23042 8632 -23008 8666
rect -22974 8632 -22940 8666
rect -22906 8632 -22872 8666
rect -22838 8632 -22804 8666
rect -22770 8632 -22736 8666
rect -22702 8632 -22668 8666
rect -22634 8632 -22600 8666
rect -22566 8632 -22532 8666
rect -22498 8632 -22464 8666
rect -22430 8632 -22396 8666
rect -22362 8632 -22328 8666
rect -22294 8632 -22260 8666
rect -22226 8632 -22192 8666
rect -22158 8632 -22124 8666
rect -22090 8632 -22056 8666
rect -22022 8632 -21988 8666
rect -21954 8632 -21920 8666
rect -21886 8632 -21852 8666
rect -21818 8632 -21784 8666
rect -21750 8632 -21716 8666
rect -21682 8632 -21648 8666
rect -21614 8632 -21580 8666
rect -21546 8632 -21512 8666
rect -21478 8632 -21444 8666
rect -21410 8632 -21376 8666
rect -21342 8632 -21308 8666
rect -21274 8632 -21240 8666
rect -21206 8632 -21172 8666
rect -21138 8632 -21104 8666
rect -21070 8632 -21036 8666
rect -21002 8632 -20968 8666
rect -20934 8632 -20900 8666
rect -20866 8632 -20832 8666
rect -20798 8632 -20764 8666
rect -20730 8632 -20696 8666
rect -20662 8632 -20628 8666
rect -20594 8632 -20560 8666
rect -20526 8632 -20492 8666
rect -20458 8632 -20424 8666
rect -20390 8632 -20356 8666
rect -20322 8632 -20288 8666
rect -20254 8632 -20220 8666
rect -20186 8632 -20152 8666
rect -20118 8632 -20084 8666
rect -20050 8632 -20016 8666
rect -19982 8632 -19948 8666
rect -19914 8632 -19880 8666
rect -19846 8632 -19812 8666
rect -19778 8632 -19744 8666
rect -19710 8632 -19676 8666
rect -19642 8632 -19608 8666
rect -19574 8632 -19540 8666
rect -19506 8632 -19472 8666
rect -19438 8632 -19404 8666
rect -19370 8632 -19336 8666
rect -19302 8632 -19268 8666
rect -19234 8632 -19200 8666
rect -19166 8632 -19132 8666
rect -19098 8632 -19064 8666
rect -19030 8632 -18996 8666
rect -18962 8632 -18928 8666
rect -18894 8632 -18860 8666
rect -18826 8632 -18792 8666
rect -18758 8632 -18724 8666
rect -18690 8632 -18656 8666
rect -18622 8632 -18588 8666
rect -18554 8632 -18520 8666
rect -18486 8632 -18452 8666
rect -18418 8632 -18384 8666
rect -18350 8632 -18316 8666
rect -18282 8632 -18248 8666
rect -18214 8632 -18180 8666
rect -18146 8632 -18112 8666
rect -18078 8632 -18044 8666
rect -18010 8632 -17976 8666
rect -17942 8632 -17908 8666
rect -17874 8632 -17840 8666
rect -17806 8632 -17772 8666
rect -17738 8632 -17704 8666
rect -17670 8632 -17636 8666
rect -17602 8632 -17568 8666
rect -17534 8632 -17500 8666
rect -17466 8632 -17432 8666
rect -17398 8632 -17364 8666
rect -17330 8632 -17296 8666
rect -17262 8632 -17228 8666
rect -17194 8632 -17160 8666
rect -17126 8632 -17092 8666
rect -17058 8632 -17024 8666
rect -16990 8632 -16956 8666
rect -16922 8632 -16888 8666
rect -16854 8632 -16820 8666
rect -16786 8632 -16752 8666
rect -16718 8632 -16684 8666
rect -16650 8632 -16616 8666
rect -16582 8632 -16548 8666
rect -16514 8632 -16480 8666
rect -16446 8632 -16412 8666
rect -16378 8632 -16344 8666
rect -16310 8632 -16276 8666
rect -16242 8632 -16208 8666
rect -16174 8632 -16140 8666
rect -16106 8632 -16072 8666
rect -16038 8632 -16004 8666
rect -15970 8632 -15936 8666
rect -15902 8632 -15868 8666
rect -15834 8632 -15800 8666
rect -15766 8632 -15732 8666
rect -15698 8632 -15664 8666
rect -15630 8632 -15596 8666
rect -15562 8632 -15528 8666
rect -15494 8632 -15460 8666
rect -15426 8632 -15392 8666
rect -15358 8632 -15324 8666
rect -15290 8632 -15256 8666
rect -15222 8632 -15188 8666
rect -15154 8632 -15120 8666
rect -15086 8632 -15052 8666
rect -15018 8632 -14984 8666
rect -14950 8632 -14916 8666
rect -14882 8632 -14848 8666
rect -14814 8632 -14780 8666
rect -14746 8632 -14712 8666
rect -14678 8632 -14644 8666
rect -14610 8632 -14576 8666
rect -14542 8632 -14508 8666
rect -14474 8632 -14440 8666
rect -14406 8632 -14372 8666
rect -14338 8632 -14304 8666
rect -14270 8632 -14236 8666
rect -14202 8632 -14168 8666
rect -14134 8632 -14100 8666
rect -14066 8632 -14032 8666
rect -13998 8632 -13964 8666
rect -13930 8632 -13896 8666
rect -13862 8632 -13828 8666
rect -13794 8632 -13760 8666
rect -13726 8632 -13692 8666
rect -13658 8632 -13624 8666
rect -13590 8632 -13360 8666
rect -26158 8466 -26124 8632
rect -26158 8398 -26124 8432
rect -26158 8330 -26124 8364
rect -26158 8262 -26124 8296
rect -26158 8194 -26124 8228
rect -26158 8126 -26124 8160
rect -26158 8058 -26124 8092
rect -26158 7990 -26124 8024
rect -26158 7922 -26124 7956
rect -26158 7854 -26124 7888
rect -26158 7786 -26124 7820
rect -26158 7718 -26124 7752
rect -26158 7650 -26124 7684
rect -26158 7582 -26124 7616
rect -26158 7514 -26124 7548
rect -26158 7446 -26124 7480
rect -26158 7378 -26124 7412
rect -26158 7310 -26124 7344
rect -26158 7242 -26124 7276
rect -26158 7174 -26124 7208
rect -26158 7106 -26124 7140
rect -26158 7038 -26124 7072
rect -26158 6970 -26124 7004
rect -26158 6902 -26124 6936
rect -26158 6834 -26124 6868
rect -26158 6766 -26124 6800
rect -26158 6698 -26124 6732
rect -26158 6630 -26124 6664
rect -26158 6562 -26124 6596
rect -26158 6494 -26124 6528
rect -26158 6426 -26124 6460
rect -26158 6358 -26124 6392
rect -26158 6290 -26124 6324
rect -26158 6222 -26124 6256
rect -26158 6154 -26124 6188
rect -26158 6086 -26124 6120
rect -26158 6018 -26124 6052
rect -26158 5950 -26124 5984
rect -26158 5882 -26124 5916
rect -26158 5814 -26124 5848
rect -26158 5746 -26124 5780
rect -26158 5678 -26124 5712
rect -26158 5610 -26124 5644
rect -26158 5542 -26124 5576
rect -26158 5325 -26124 5508
rect -13394 8466 -13360 8632
rect -13394 8398 -13360 8432
rect -13394 8330 -13360 8364
rect -13394 8262 -13360 8296
rect -13394 8194 -13360 8228
rect -13394 8126 -13360 8160
rect -13394 8058 -13360 8092
rect -13394 7990 -13360 8024
rect -13394 7922 -13360 7956
rect -13394 7854 -13360 7888
rect -13394 7786 -13360 7820
rect -13394 7718 -13360 7752
rect -13394 7650 -13360 7684
rect -13394 7582 -13360 7616
rect -13394 7514 -13360 7548
rect -13394 7446 -13360 7480
rect -13394 7378 -13360 7412
rect -13394 7310 -13360 7344
rect -13394 7242 -13360 7276
rect -13394 7174 -13360 7208
rect -13394 7106 -13360 7140
rect -13394 7038 -13360 7072
rect -13394 6970 -13360 7004
rect -13394 6902 -13360 6936
rect -13394 6834 -13360 6868
rect -13394 6766 -13360 6800
rect -13394 6698 -13360 6732
rect -13394 6630 -13360 6664
rect -13394 6562 -13360 6596
rect -13394 6494 -13360 6528
rect -13394 6426 -13360 6460
rect -13394 6358 -13360 6392
rect -13394 6290 -13360 6324
rect -13394 6222 -13360 6256
rect -13394 6154 -13360 6188
rect -13394 6086 -13360 6120
rect -13394 6018 -13360 6052
rect -13394 5950 -13360 5984
rect -13394 5882 -13360 5916
rect -13394 5814 -13360 5848
rect -13394 5746 -13360 5780
rect -13394 5678 -13360 5712
rect -13394 5610 -13360 5644
rect -13394 5542 -13360 5576
rect -13394 5325 -13360 5508
rect -26158 5291 -25958 5325
rect -25924 5291 -25890 5325
rect -25856 5291 -25822 5325
rect -25788 5291 -25754 5325
rect -25720 5291 -25686 5325
rect -25652 5291 -25618 5325
rect -25584 5291 -25550 5325
rect -25516 5291 -25482 5325
rect -25448 5291 -25414 5325
rect -25380 5291 -25346 5325
rect -25312 5291 -25278 5325
rect -25244 5291 -25210 5325
rect -25176 5291 -25142 5325
rect -25108 5291 -25074 5325
rect -25040 5291 -25006 5325
rect -24972 5291 -24938 5325
rect -24904 5291 -24870 5325
rect -24836 5291 -24802 5325
rect -24768 5291 -24734 5325
rect -24700 5291 -24666 5325
rect -24632 5291 -24598 5325
rect -24564 5291 -24530 5325
rect -24496 5291 -24462 5325
rect -24428 5291 -24394 5325
rect -24360 5291 -24326 5325
rect -24292 5291 -24258 5325
rect -24224 5291 -24190 5325
rect -24156 5291 -24122 5325
rect -24088 5291 -24054 5325
rect -24020 5291 -23986 5325
rect -23952 5291 -23918 5325
rect -23884 5291 -23850 5325
rect -23816 5291 -23782 5325
rect -23748 5291 -23714 5325
rect -23680 5291 -23646 5325
rect -23612 5291 -23578 5325
rect -23544 5291 -23510 5325
rect -23476 5291 -23442 5325
rect -23408 5291 -23374 5325
rect -23340 5291 -23306 5325
rect -23272 5291 -23238 5325
rect -23204 5291 -23170 5325
rect -23136 5291 -23102 5325
rect -23068 5291 -23034 5325
rect -23000 5291 -22966 5325
rect -22932 5291 -22898 5325
rect -22864 5291 -22830 5325
rect -22796 5291 -22762 5325
rect -22728 5291 -22694 5325
rect -22660 5291 -22626 5325
rect -22592 5291 -22558 5325
rect -22524 5291 -22490 5325
rect -22456 5291 -22422 5325
rect -22388 5291 -22354 5325
rect -22320 5291 -22286 5325
rect -22252 5291 -22218 5325
rect -22184 5291 -22150 5325
rect -22116 5291 -22082 5325
rect -22048 5291 -22014 5325
rect -21980 5291 -21946 5325
rect -21912 5291 -21878 5325
rect -21844 5291 -21810 5325
rect -21776 5291 -21742 5325
rect -21708 5291 -21674 5325
rect -21640 5291 -21606 5325
rect -21572 5291 -21538 5325
rect -21504 5291 -21470 5325
rect -21436 5291 -21402 5325
rect -21368 5291 -21334 5325
rect -21300 5291 -21266 5325
rect -21232 5291 -21198 5325
rect -21164 5291 -21130 5325
rect -21096 5291 -21062 5325
rect -21028 5291 -20994 5325
rect -20960 5291 -20926 5325
rect -20892 5291 -20858 5325
rect -20824 5291 -20790 5325
rect -20756 5291 -20722 5325
rect -20688 5291 -20654 5325
rect -20620 5291 -20586 5325
rect -20552 5291 -20518 5325
rect -20484 5291 -20450 5325
rect -20416 5291 -20382 5325
rect -20348 5291 -20314 5325
rect -20280 5291 -20246 5325
rect -20212 5291 -20178 5325
rect -20144 5291 -20110 5325
rect -20076 5291 -20042 5325
rect -20008 5291 -19974 5325
rect -19940 5291 -19906 5325
rect -19872 5291 -19838 5325
rect -19804 5291 -19770 5325
rect -19736 5291 -19702 5325
rect -19668 5291 -19634 5325
rect -19600 5291 -19566 5325
rect -19532 5291 -19498 5325
rect -19464 5291 -19430 5325
rect -19396 5291 -19362 5325
rect -19328 5291 -19294 5325
rect -19260 5291 -19226 5325
rect -19192 5291 -19158 5325
rect -19124 5291 -19090 5325
rect -19056 5291 -19022 5325
rect -18988 5291 -18954 5325
rect -18920 5291 -18886 5325
rect -18852 5291 -18818 5325
rect -18784 5291 -18750 5325
rect -18716 5291 -18682 5325
rect -18648 5291 -18614 5325
rect -18580 5291 -18546 5325
rect -18512 5291 -18478 5325
rect -18444 5291 -18410 5325
rect -18376 5291 -18342 5325
rect -18308 5291 -18274 5325
rect -18240 5291 -18206 5325
rect -18172 5291 -18138 5325
rect -18104 5291 -18070 5325
rect -18036 5291 -18002 5325
rect -17968 5291 -17934 5325
rect -17900 5291 -17866 5325
rect -17832 5291 -17798 5325
rect -17764 5291 -17730 5325
rect -17696 5291 -17662 5325
rect -17628 5291 -17594 5325
rect -17560 5291 -17526 5325
rect -17492 5291 -17458 5325
rect -17424 5291 -17390 5325
rect -17356 5291 -17322 5325
rect -17288 5291 -17254 5325
rect -17220 5291 -17186 5325
rect -17152 5291 -17118 5325
rect -17084 5291 -17050 5325
rect -17016 5291 -16982 5325
rect -16948 5291 -16914 5325
rect -16880 5291 -16846 5325
rect -16812 5291 -16778 5325
rect -16744 5291 -16710 5325
rect -16676 5291 -16642 5325
rect -16608 5291 -16574 5325
rect -16540 5291 -16506 5325
rect -16472 5291 -16438 5325
rect -16404 5291 -16370 5325
rect -16336 5291 -16302 5325
rect -16268 5291 -16234 5325
rect -16200 5291 -16166 5325
rect -16132 5291 -16098 5325
rect -16064 5291 -16030 5325
rect -15996 5291 -15962 5325
rect -15928 5291 -15894 5325
rect -15860 5291 -15826 5325
rect -15792 5291 -15758 5325
rect -15724 5291 -15690 5325
rect -15656 5291 -15622 5325
rect -15588 5291 -15554 5325
rect -15520 5291 -15486 5325
rect -15452 5291 -15418 5325
rect -15384 5291 -15350 5325
rect -15316 5291 -15282 5325
rect -15248 5291 -15214 5325
rect -15180 5291 -15146 5325
rect -15112 5291 -15078 5325
rect -15044 5291 -15010 5325
rect -14976 5291 -14942 5325
rect -14908 5291 -14874 5325
rect -14840 5291 -14806 5325
rect -14772 5291 -14738 5325
rect -14704 5291 -14670 5325
rect -14636 5291 -14602 5325
rect -14568 5291 -14534 5325
rect -14500 5291 -14466 5325
rect -14432 5291 -14398 5325
rect -14364 5291 -14330 5325
rect -14296 5291 -14262 5325
rect -14228 5291 -14194 5325
rect -14160 5291 -14126 5325
rect -14092 5291 -14058 5325
rect -14024 5291 -13990 5325
rect -13956 5291 -13922 5325
rect -13888 5291 -13854 5325
rect -13820 5291 -13786 5325
rect -13752 5291 -13718 5325
rect -13684 5291 -13650 5325
rect -13616 5291 -13360 5325
<< properties >>
string path -130.915 43.245 -66.885 43.245 -66.885 26.540 -130.705 26.540 -130.705 43.245 
<< end >>
