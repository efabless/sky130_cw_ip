magic
tech sky130A
magscale 1 2
timestamp 1715010268
<< nwell >>
rect -314 2942 3090 3110
rect -314 -126 -146 2942
rect 2922 -126 3090 2942
rect -314 -294 3090 -126
<< nsubdiff >>
rect -247 3009 -143 3043
rect -109 3009 -75 3043
rect -41 3009 -7 3043
rect 27 3009 61 3043
rect 95 3009 129 3043
rect 163 3009 197 3043
rect 231 3009 265 3043
rect 299 3009 333 3043
rect 367 3009 401 3043
rect 435 3009 469 3043
rect 503 3009 537 3043
rect 571 3009 605 3043
rect 639 3009 673 3043
rect 707 3009 741 3043
rect 775 3009 809 3043
rect 843 3009 877 3043
rect 911 3009 945 3043
rect 979 3009 1013 3043
rect 1047 3009 1081 3043
rect 1115 3009 1149 3043
rect 1183 3009 1217 3043
rect 1251 3009 1285 3043
rect 1319 3009 1353 3043
rect 1387 3009 1421 3043
rect 1455 3009 1489 3043
rect 1523 3009 1557 3043
rect 1591 3009 1625 3043
rect 1659 3009 1693 3043
rect 1727 3009 1761 3043
rect 1795 3009 1829 3043
rect 1863 3009 1897 3043
rect 1931 3009 1965 3043
rect 1999 3009 2033 3043
rect 2067 3009 2101 3043
rect 2135 3009 2169 3043
rect 2203 3009 2237 3043
rect 2271 3009 2305 3043
rect 2339 3009 2373 3043
rect 2407 3009 2441 3043
rect 2475 3009 2509 3043
rect 2543 3009 2577 3043
rect 2611 3009 2645 3043
rect 2679 3009 2713 3043
rect 2747 3009 2781 3043
rect 2815 3009 2849 3043
rect 2883 3009 3023 3043
rect -247 2903 -213 3009
rect -247 2835 -213 2869
rect -247 2767 -213 2801
rect -247 2699 -213 2733
rect -247 2631 -213 2665
rect -247 2563 -213 2597
rect -247 2495 -213 2529
rect -247 2427 -213 2461
rect -247 2359 -213 2393
rect -247 2291 -213 2325
rect -247 2223 -213 2257
rect -247 2155 -213 2189
rect -247 2087 -213 2121
rect -247 2019 -213 2053
rect -247 1951 -213 1985
rect -247 1883 -213 1917
rect -247 1815 -213 1849
rect -247 1747 -213 1781
rect -247 1679 -213 1713
rect -247 1611 -213 1645
rect -247 1543 -213 1577
rect -247 1475 -213 1509
rect -247 1407 -213 1441
rect -247 1339 -213 1373
rect -247 1271 -213 1305
rect -247 1203 -213 1237
rect -247 1135 -213 1169
rect -247 1067 -213 1101
rect -247 999 -213 1033
rect -247 931 -213 965
rect -247 863 -213 897
rect -247 795 -213 829
rect -247 727 -213 761
rect -247 659 -213 693
rect -247 591 -213 625
rect -247 523 -213 557
rect -247 455 -213 489
rect -247 387 -213 421
rect -247 319 -213 353
rect -247 251 -213 285
rect -247 183 -213 217
rect -247 115 -213 149
rect -247 47 -213 81
rect -247 -21 -213 13
rect -247 -193 -213 -55
rect 2989 2903 3023 3009
rect 2989 2835 3023 2869
rect 2989 2767 3023 2801
rect 2989 2699 3023 2733
rect 2989 2631 3023 2665
rect 2989 2563 3023 2597
rect 2989 2495 3023 2529
rect 2989 2427 3023 2461
rect 2989 2359 3023 2393
rect 2989 2291 3023 2325
rect 2989 2223 3023 2257
rect 2989 2155 3023 2189
rect 2989 2087 3023 2121
rect 2989 2019 3023 2053
rect 2989 1951 3023 1985
rect 2989 1883 3023 1917
rect 2989 1815 3023 1849
rect 2989 1747 3023 1781
rect 2989 1679 3023 1713
rect 2989 1611 3023 1645
rect 2989 1543 3023 1577
rect 2989 1475 3023 1509
rect 2989 1407 3023 1441
rect 2989 1339 3023 1373
rect 2989 1271 3023 1305
rect 2989 1203 3023 1237
rect 2989 1135 3023 1169
rect 2989 1067 3023 1101
rect 2989 999 3023 1033
rect 2989 931 3023 965
rect 2989 863 3023 897
rect 2989 795 3023 829
rect 2989 727 3023 761
rect 2989 659 3023 693
rect 2989 591 3023 625
rect 2989 523 3023 557
rect 2989 455 3023 489
rect 2989 387 3023 421
rect 2989 319 3023 353
rect 2989 251 3023 285
rect 2989 183 3023 217
rect 2989 115 3023 149
rect 2989 47 3023 81
rect 2989 -21 3023 13
rect 2989 -193 3023 -55
rect -247 -227 -75 -193
rect -41 -227 -7 -193
rect 27 -227 61 -193
rect 95 -227 129 -193
rect 163 -227 197 -193
rect 231 -227 265 -193
rect 299 -227 333 -193
rect 367 -227 401 -193
rect 435 -227 469 -193
rect 503 -227 537 -193
rect 571 -227 605 -193
rect 639 -227 673 -193
rect 707 -227 741 -193
rect 775 -227 809 -193
rect 843 -227 877 -193
rect 911 -227 945 -193
rect 979 -227 1013 -193
rect 1047 -227 1081 -193
rect 1115 -227 1149 -193
rect 1183 -227 1217 -193
rect 1251 -227 1285 -193
rect 1319 -227 1353 -193
rect 1387 -227 1421 -193
rect 1455 -227 1489 -193
rect 1523 -227 1557 -193
rect 1591 -227 1625 -193
rect 1659 -227 1693 -193
rect 1727 -227 1761 -193
rect 1795 -227 1829 -193
rect 1863 -227 1897 -193
rect 1931 -227 1965 -193
rect 1999 -227 2033 -193
rect 2067 -227 2101 -193
rect 2135 -227 2169 -193
rect 2203 -227 2237 -193
rect 2271 -227 2305 -193
rect 2339 -227 2373 -193
rect 2407 -227 2441 -193
rect 2475 -227 2509 -193
rect 2543 -227 2577 -193
rect 2611 -227 2645 -193
rect 2679 -227 2713 -193
rect 2747 -227 2781 -193
rect 2815 -227 2849 -193
rect 2883 -227 3023 -193
<< nsubdiffcont >>
rect -143 3009 -109 3043
rect -75 3009 -41 3043
rect -7 3009 27 3043
rect 61 3009 95 3043
rect 129 3009 163 3043
rect 197 3009 231 3043
rect 265 3009 299 3043
rect 333 3009 367 3043
rect 401 3009 435 3043
rect 469 3009 503 3043
rect 537 3009 571 3043
rect 605 3009 639 3043
rect 673 3009 707 3043
rect 741 3009 775 3043
rect 809 3009 843 3043
rect 877 3009 911 3043
rect 945 3009 979 3043
rect 1013 3009 1047 3043
rect 1081 3009 1115 3043
rect 1149 3009 1183 3043
rect 1217 3009 1251 3043
rect 1285 3009 1319 3043
rect 1353 3009 1387 3043
rect 1421 3009 1455 3043
rect 1489 3009 1523 3043
rect 1557 3009 1591 3043
rect 1625 3009 1659 3043
rect 1693 3009 1727 3043
rect 1761 3009 1795 3043
rect 1829 3009 1863 3043
rect 1897 3009 1931 3043
rect 1965 3009 1999 3043
rect 2033 3009 2067 3043
rect 2101 3009 2135 3043
rect 2169 3009 2203 3043
rect 2237 3009 2271 3043
rect 2305 3009 2339 3043
rect 2373 3009 2407 3043
rect 2441 3009 2475 3043
rect 2509 3009 2543 3043
rect 2577 3009 2611 3043
rect 2645 3009 2679 3043
rect 2713 3009 2747 3043
rect 2781 3009 2815 3043
rect 2849 3009 2883 3043
rect -247 2869 -213 2903
rect -247 2801 -213 2835
rect -247 2733 -213 2767
rect -247 2665 -213 2699
rect -247 2597 -213 2631
rect -247 2529 -213 2563
rect -247 2461 -213 2495
rect -247 2393 -213 2427
rect -247 2325 -213 2359
rect -247 2257 -213 2291
rect -247 2189 -213 2223
rect -247 2121 -213 2155
rect -247 2053 -213 2087
rect -247 1985 -213 2019
rect -247 1917 -213 1951
rect -247 1849 -213 1883
rect -247 1781 -213 1815
rect -247 1713 -213 1747
rect -247 1645 -213 1679
rect -247 1577 -213 1611
rect -247 1509 -213 1543
rect -247 1441 -213 1475
rect -247 1373 -213 1407
rect -247 1305 -213 1339
rect -247 1237 -213 1271
rect -247 1169 -213 1203
rect -247 1101 -213 1135
rect -247 1033 -213 1067
rect -247 965 -213 999
rect -247 897 -213 931
rect -247 829 -213 863
rect -247 761 -213 795
rect -247 693 -213 727
rect -247 625 -213 659
rect -247 557 -213 591
rect -247 489 -213 523
rect -247 421 -213 455
rect -247 353 -213 387
rect -247 285 -213 319
rect -247 217 -213 251
rect -247 149 -213 183
rect -247 81 -213 115
rect -247 13 -213 47
rect -247 -55 -213 -21
rect 2989 2869 3023 2903
rect 2989 2801 3023 2835
rect 2989 2733 3023 2767
rect 2989 2665 3023 2699
rect 2989 2597 3023 2631
rect 2989 2529 3023 2563
rect 2989 2461 3023 2495
rect 2989 2393 3023 2427
rect 2989 2325 3023 2359
rect 2989 2257 3023 2291
rect 2989 2189 3023 2223
rect 2989 2121 3023 2155
rect 2989 2053 3023 2087
rect 2989 1985 3023 2019
rect 2989 1917 3023 1951
rect 2989 1849 3023 1883
rect 2989 1781 3023 1815
rect 2989 1713 3023 1747
rect 2989 1645 3023 1679
rect 2989 1577 3023 1611
rect 2989 1509 3023 1543
rect 2989 1441 3023 1475
rect 2989 1373 3023 1407
rect 2989 1305 3023 1339
rect 2989 1237 3023 1271
rect 2989 1169 3023 1203
rect 2989 1101 3023 1135
rect 2989 1033 3023 1067
rect 2989 965 3023 999
rect 2989 897 3023 931
rect 2989 829 3023 863
rect 2989 761 3023 795
rect 2989 693 3023 727
rect 2989 625 3023 659
rect 2989 557 3023 591
rect 2989 489 3023 523
rect 2989 421 3023 455
rect 2989 353 3023 387
rect 2989 285 3023 319
rect 2989 217 3023 251
rect 2989 149 3023 183
rect 2989 81 3023 115
rect 2989 13 3023 47
rect 2989 -55 3023 -21
rect -75 -227 -41 -193
rect -7 -227 27 -193
rect 61 -227 95 -193
rect 129 -227 163 -193
rect 197 -227 231 -193
rect 265 -227 299 -193
rect 333 -227 367 -193
rect 401 -227 435 -193
rect 469 -227 503 -193
rect 537 -227 571 -193
rect 605 -227 639 -193
rect 673 -227 707 -193
rect 741 -227 775 -193
rect 809 -227 843 -193
rect 877 -227 911 -193
rect 945 -227 979 -193
rect 1013 -227 1047 -193
rect 1081 -227 1115 -193
rect 1149 -227 1183 -193
rect 1217 -227 1251 -193
rect 1285 -227 1319 -193
rect 1353 -227 1387 -193
rect 1421 -227 1455 -193
rect 1489 -227 1523 -193
rect 1557 -227 1591 -193
rect 1625 -227 1659 -193
rect 1693 -227 1727 -193
rect 1761 -227 1795 -193
rect 1829 -227 1863 -193
rect 1897 -227 1931 -193
rect 1965 -227 1999 -193
rect 2033 -227 2067 -193
rect 2101 -227 2135 -193
rect 2169 -227 2203 -193
rect 2237 -227 2271 -193
rect 2305 -227 2339 -193
rect 2373 -227 2407 -193
rect 2441 -227 2475 -193
rect 2509 -227 2543 -193
rect 2577 -227 2611 -193
rect 2645 -227 2679 -193
rect 2713 -227 2747 -193
rect 2781 -227 2815 -193
rect 2849 -227 2883 -193
<< locali >>
rect -247 3009 -143 3043
rect -109 3009 -75 3043
rect -41 3009 -7 3043
rect 27 3009 61 3043
rect 95 3009 129 3043
rect 163 3009 197 3043
rect 231 3009 265 3043
rect 299 3009 333 3043
rect 367 3009 401 3043
rect 435 3009 469 3043
rect 503 3009 537 3043
rect 571 3009 605 3043
rect 639 3009 673 3043
rect 707 3009 741 3043
rect 775 3009 809 3043
rect 843 3009 877 3043
rect 911 3009 945 3043
rect 979 3009 1013 3043
rect 1047 3009 1081 3043
rect 1115 3009 1149 3043
rect 1183 3009 1217 3043
rect 1251 3009 1285 3043
rect 1319 3009 1353 3043
rect 1387 3009 1421 3043
rect 1455 3009 1489 3043
rect 1523 3009 1557 3043
rect 1591 3009 1625 3043
rect 1659 3009 1693 3043
rect 1727 3009 1761 3043
rect 1795 3009 1829 3043
rect 1863 3009 1897 3043
rect 1931 3009 1965 3043
rect 1999 3009 2033 3043
rect 2067 3009 2101 3043
rect 2135 3009 2169 3043
rect 2203 3009 2237 3043
rect 2271 3009 2305 3043
rect 2339 3009 2373 3043
rect 2407 3009 2441 3043
rect 2475 3009 2509 3043
rect 2543 3009 2577 3043
rect 2611 3009 2645 3043
rect 2679 3009 2713 3043
rect 2747 3009 2781 3043
rect 2815 3009 2849 3043
rect 2883 3009 3023 3043
rect -247 2903 -213 3009
rect -247 2835 -213 2869
rect -247 2767 -213 2801
rect -247 2699 -213 2733
rect -247 2631 -213 2665
rect -247 2563 -213 2597
rect -247 2495 -213 2529
rect -247 2427 -213 2461
rect -247 2359 -213 2393
rect -247 2291 -213 2325
rect -247 2223 -213 2257
rect -247 2155 -213 2189
rect -247 2087 -213 2121
rect -247 2019 -213 2053
rect -247 1951 -213 1985
rect -247 1883 -213 1917
rect -247 1815 -213 1849
rect -247 1747 -213 1781
rect -247 1679 -213 1713
rect -247 1611 -213 1645
rect -247 1543 -213 1577
rect -247 1475 -213 1509
rect -247 1407 -213 1441
rect -247 1339 -213 1373
rect -247 1271 -213 1305
rect -247 1203 -213 1237
rect -247 1135 -213 1169
rect -247 1067 -213 1101
rect -247 999 -213 1033
rect -247 931 -213 965
rect -247 863 -213 897
rect -247 795 -213 829
rect -247 727 -213 761
rect -247 659 -213 693
rect -247 591 -213 625
rect -247 523 -213 557
rect -247 455 -213 489
rect -247 387 -213 421
rect -247 319 -213 353
rect -247 251 -213 285
rect -247 183 -213 217
rect -247 115 -213 149
rect -247 47 -213 81
rect -247 -21 -213 13
rect -247 -193 -213 -55
rect 2989 2903 3023 3009
rect 2989 2835 3023 2869
rect 2989 2767 3023 2801
rect 2989 2699 3023 2733
rect 2989 2631 3023 2665
rect 2989 2563 3023 2597
rect 2989 2495 3023 2529
rect 2989 2427 3023 2461
rect 2989 2359 3023 2393
rect 2989 2291 3023 2325
rect 2989 2223 3023 2257
rect 2989 2155 3023 2189
rect 2989 2087 3023 2121
rect 2989 2019 3023 2053
rect 2989 1951 3023 1985
rect 2989 1883 3023 1917
rect 2989 1815 3023 1849
rect 2989 1747 3023 1781
rect 2989 1679 3023 1713
rect 2989 1611 3023 1645
rect 2989 1543 3023 1577
rect 2989 1475 3023 1509
rect 2989 1407 3023 1441
rect 2989 1339 3023 1373
rect 2989 1271 3023 1305
rect 2989 1203 3023 1237
rect 2989 1135 3023 1169
rect 2989 1067 3023 1101
rect 2989 999 3023 1033
rect 2989 931 3023 965
rect 2989 863 3023 897
rect 2989 795 3023 829
rect 2989 727 3023 761
rect 2989 659 3023 693
rect 2989 591 3023 625
rect 2989 523 3023 557
rect 2989 455 3023 489
rect 2989 387 3023 421
rect 2989 319 3023 353
rect 2989 251 3023 285
rect 2989 183 3023 217
rect 2989 115 3023 149
rect 2989 47 3023 81
rect 2989 -21 3023 13
rect 2989 -193 3023 -55
rect -247 -227 -75 -193
rect -41 -227 -7 -193
rect 27 -227 61 -193
rect 95 -227 129 -193
rect 163 -227 197 -193
rect 231 -227 265 -193
rect 299 -227 333 -193
rect 367 -227 401 -193
rect 435 -227 469 -193
rect 503 -227 537 -193
rect 571 -227 605 -193
rect 639 -227 673 -193
rect 707 -227 741 -193
rect 775 -227 809 -193
rect 843 -227 877 -193
rect 911 -227 945 -193
rect 979 -227 1013 -193
rect 1047 -227 1081 -193
rect 1115 -227 1149 -193
rect 1183 -227 1217 -193
rect 1251 -227 1285 -193
rect 1319 -227 1353 -193
rect 1387 -227 1421 -193
rect 1455 -227 1489 -193
rect 1523 -227 1557 -193
rect 1591 -227 1625 -193
rect 1659 -227 1693 -193
rect 1727 -227 1761 -193
rect 1795 -227 1829 -193
rect 1863 -227 1897 -193
rect 1931 -227 1965 -193
rect 1999 -227 2033 -193
rect 2067 -227 2101 -193
rect 2135 -227 2169 -193
rect 2203 -227 2237 -193
rect 2271 -227 2305 -193
rect 2339 -227 2373 -193
rect 2407 -227 2441 -193
rect 2475 -227 2509 -193
rect 2543 -227 2577 -193
rect 2611 -227 2645 -193
rect 2679 -227 2713 -193
rect 2747 -227 2781 -193
rect 2815 -227 2849 -193
rect 2883 -227 3023 -193
<< properties >>
string path -7.075 75.650 75.150 75.650 75.150 -5.250 -5.750 -5.250 -5.750 77.750 
<< end >>
