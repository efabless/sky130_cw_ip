magic
tech sky130A
magscale 1 2
timestamp 1715625863
<< metal3 >>
rect -1150 1072 1149 1100
rect -1150 1008 1065 1072
rect 1129 1008 1149 1072
rect -1150 992 1149 1008
rect -1150 928 1065 992
rect 1129 928 1149 992
rect -1150 912 1149 928
rect -1150 848 1065 912
rect 1129 848 1149 912
rect -1150 832 1149 848
rect -1150 768 1065 832
rect 1129 768 1149 832
rect -1150 752 1149 768
rect -1150 688 1065 752
rect 1129 688 1149 752
rect -1150 672 1149 688
rect -1150 608 1065 672
rect 1129 608 1149 672
rect -1150 592 1149 608
rect -1150 528 1065 592
rect 1129 528 1149 592
rect -1150 512 1149 528
rect -1150 448 1065 512
rect 1129 448 1149 512
rect -1150 432 1149 448
rect -1150 368 1065 432
rect 1129 368 1149 432
rect -1150 352 1149 368
rect -1150 288 1065 352
rect 1129 288 1149 352
rect -1150 272 1149 288
rect -1150 208 1065 272
rect 1129 208 1149 272
rect -1150 192 1149 208
rect -1150 128 1065 192
rect 1129 128 1149 192
rect -1150 112 1149 128
rect -1150 48 1065 112
rect 1129 48 1149 112
rect -1150 32 1149 48
rect -1150 -32 1065 32
rect 1129 -32 1149 32
rect -1150 -48 1149 -32
rect -1150 -112 1065 -48
rect 1129 -112 1149 -48
rect -1150 -128 1149 -112
rect -1150 -192 1065 -128
rect 1129 -192 1149 -128
rect -1150 -208 1149 -192
rect -1150 -272 1065 -208
rect 1129 -272 1149 -208
rect -1150 -288 1149 -272
rect -1150 -352 1065 -288
rect 1129 -352 1149 -288
rect -1150 -368 1149 -352
rect -1150 -432 1065 -368
rect 1129 -432 1149 -368
rect -1150 -448 1149 -432
rect -1150 -512 1065 -448
rect 1129 -512 1149 -448
rect -1150 -528 1149 -512
rect -1150 -592 1065 -528
rect 1129 -592 1149 -528
rect -1150 -608 1149 -592
rect -1150 -672 1065 -608
rect 1129 -672 1149 -608
rect -1150 -688 1149 -672
rect -1150 -752 1065 -688
rect 1129 -752 1149 -688
rect -1150 -768 1149 -752
rect -1150 -832 1065 -768
rect 1129 -832 1149 -768
rect -1150 -848 1149 -832
rect -1150 -912 1065 -848
rect 1129 -912 1149 -848
rect -1150 -928 1149 -912
rect -1150 -992 1065 -928
rect 1129 -992 1149 -928
rect -1150 -1008 1149 -992
rect -1150 -1072 1065 -1008
rect 1129 -1072 1149 -1008
rect -1150 -1100 1149 -1072
<< via3 >>
rect 1065 1008 1129 1072
rect 1065 928 1129 992
rect 1065 848 1129 912
rect 1065 768 1129 832
rect 1065 688 1129 752
rect 1065 608 1129 672
rect 1065 528 1129 592
rect 1065 448 1129 512
rect 1065 368 1129 432
rect 1065 288 1129 352
rect 1065 208 1129 272
rect 1065 128 1129 192
rect 1065 48 1129 112
rect 1065 -32 1129 32
rect 1065 -112 1129 -48
rect 1065 -192 1129 -128
rect 1065 -272 1129 -208
rect 1065 -352 1129 -288
rect 1065 -432 1129 -368
rect 1065 -512 1129 -448
rect 1065 -592 1129 -528
rect 1065 -672 1129 -608
rect 1065 -752 1129 -688
rect 1065 -832 1129 -768
rect 1065 -912 1129 -848
rect 1065 -992 1129 -928
rect 1065 -1072 1129 -1008
<< mimcap >>
rect -1050 952 950 1000
rect -1050 -952 -1002 952
rect 902 -952 950 952
rect -1050 -1000 950 -952
<< mimcapcontact >>
rect -1002 -952 902 952
<< metal4 >>
rect 1049 1072 1145 1088
rect 1049 1008 1065 1072
rect 1129 1008 1145 1072
rect 1049 992 1145 1008
rect -1011 952 911 961
rect -1011 -952 -1002 952
rect 902 -952 911 952
rect -1011 -961 911 -952
rect 1049 928 1065 992
rect 1129 928 1145 992
rect 1049 912 1145 928
rect 1049 848 1065 912
rect 1129 848 1145 912
rect 1049 832 1145 848
rect 1049 768 1065 832
rect 1129 768 1145 832
rect 1049 752 1145 768
rect 1049 688 1065 752
rect 1129 688 1145 752
rect 1049 672 1145 688
rect 1049 608 1065 672
rect 1129 608 1145 672
rect 1049 592 1145 608
rect 1049 528 1065 592
rect 1129 528 1145 592
rect 1049 512 1145 528
rect 1049 448 1065 512
rect 1129 448 1145 512
rect 1049 432 1145 448
rect 1049 368 1065 432
rect 1129 368 1145 432
rect 1049 352 1145 368
rect 1049 288 1065 352
rect 1129 288 1145 352
rect 1049 272 1145 288
rect 1049 208 1065 272
rect 1129 208 1145 272
rect 1049 192 1145 208
rect 1049 128 1065 192
rect 1129 128 1145 192
rect 1049 112 1145 128
rect 1049 48 1065 112
rect 1129 48 1145 112
rect 1049 32 1145 48
rect 1049 -32 1065 32
rect 1129 -32 1145 32
rect 1049 -48 1145 -32
rect 1049 -112 1065 -48
rect 1129 -112 1145 -48
rect 1049 -128 1145 -112
rect 1049 -192 1065 -128
rect 1129 -192 1145 -128
rect 1049 -208 1145 -192
rect 1049 -272 1065 -208
rect 1129 -272 1145 -208
rect 1049 -288 1145 -272
rect 1049 -352 1065 -288
rect 1129 -352 1145 -288
rect 1049 -368 1145 -352
rect 1049 -432 1065 -368
rect 1129 -432 1145 -368
rect 1049 -448 1145 -432
rect 1049 -512 1065 -448
rect 1129 -512 1145 -448
rect 1049 -528 1145 -512
rect 1049 -592 1065 -528
rect 1129 -592 1145 -528
rect 1049 -608 1145 -592
rect 1049 -672 1065 -608
rect 1129 -672 1145 -608
rect 1049 -688 1145 -672
rect 1049 -752 1065 -688
rect 1129 -752 1145 -688
rect 1049 -768 1145 -752
rect 1049 -832 1065 -768
rect 1129 -832 1145 -768
rect 1049 -848 1145 -832
rect 1049 -912 1065 -848
rect 1129 -912 1145 -848
rect 1049 -928 1145 -912
rect 1049 -992 1065 -928
rect 1129 -992 1145 -928
rect 1049 -1008 1145 -992
rect 1049 -1072 1065 -1008
rect 1129 -1072 1145 -1008
rect 1049 -1088 1145 -1072
<< properties >>
string FIXED_BBOX -1150 -1100 1050 1100
<< end >>
