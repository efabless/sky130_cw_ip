magic
tech sky130A
magscale 1 2
timestamp 1715010268
<< pwell >>
rect -184 -157 184 95
<< nmoslvt >>
rect -100 -131 100 69
<< ndiff >>
rect -158 54 -100 69
rect -158 20 -146 54
rect -112 20 -100 54
rect -158 -14 -100 20
rect -158 -48 -146 -14
rect -112 -48 -100 -14
rect -158 -82 -100 -48
rect -158 -116 -146 -82
rect -112 -116 -100 -82
rect -158 -131 -100 -116
rect 100 54 158 69
rect 100 20 112 54
rect 146 20 158 54
rect 100 -14 158 20
rect 100 -48 112 -14
rect 146 -48 158 -14
rect 100 -82 158 -48
rect 100 -116 112 -82
rect 146 -116 158 -82
rect 100 -131 158 -116
<< ndiffc >>
rect -146 20 -112 54
rect -146 -48 -112 -14
rect -146 -116 -112 -82
rect 112 20 146 54
rect 112 -48 146 -14
rect 112 -116 146 -82
<< poly >>
rect -100 141 100 157
rect -100 107 -51 141
rect -17 107 17 141
rect 51 107 100 141
rect -100 69 100 107
rect -100 -157 100 -131
<< polycont >>
rect -51 107 -17 141
rect 17 107 51 141
<< locali >>
rect -100 107 -53 141
rect -17 107 17 141
rect 53 107 100 141
rect -146 54 -112 73
rect -146 -14 -112 -12
rect -146 -50 -112 -48
rect -146 -135 -112 -116
rect 112 54 146 73
rect 112 -14 146 -12
rect 112 -50 146 -48
rect 112 -135 146 -116
<< viali >>
rect -53 107 -51 141
rect -51 107 -19 141
rect 19 107 51 141
rect 51 107 53 141
rect -146 20 -112 22
rect -146 -12 -112 20
rect -146 -82 -112 -50
rect -146 -84 -112 -82
rect 112 20 146 22
rect 112 -12 146 20
rect 112 -82 146 -50
rect 112 -84 146 -82
<< metal1 >>
rect -96 141 96 147
rect -96 107 -53 141
rect -19 107 19 141
rect 53 107 96 141
rect -96 101 96 107
rect -152 22 -106 69
rect -152 -12 -146 22
rect -112 -12 -106 22
rect -152 -50 -106 -12
rect -152 -84 -146 -50
rect -112 -84 -106 -50
rect -152 -131 -106 -84
rect 106 22 152 69
rect 106 -12 112 22
rect 146 -12 152 22
rect 106 -50 152 -12
rect 106 -84 112 -50
rect 146 -84 152 -50
rect 106 -131 152 -84
<< end >>
