magic
tech sky130A
magscale 1 2
timestamp 1715625863
<< error_p >>
rect -194 -498 194 464
<< nwell >>
rect -194 -498 194 464
<< pmoslvt >>
rect -100 -436 100 364
<< pdiff >>
rect -158 321 -100 364
rect -158 287 -146 321
rect -112 287 -100 321
rect -158 253 -100 287
rect -158 219 -146 253
rect -112 219 -100 253
rect -158 185 -100 219
rect -158 151 -146 185
rect -112 151 -100 185
rect -158 117 -100 151
rect -158 83 -146 117
rect -112 83 -100 117
rect -158 49 -100 83
rect -158 15 -146 49
rect -112 15 -100 49
rect -158 -19 -100 15
rect -158 -53 -146 -19
rect -112 -53 -100 -19
rect -158 -87 -100 -53
rect -158 -121 -146 -87
rect -112 -121 -100 -87
rect -158 -155 -100 -121
rect -158 -189 -146 -155
rect -112 -189 -100 -155
rect -158 -223 -100 -189
rect -158 -257 -146 -223
rect -112 -257 -100 -223
rect -158 -291 -100 -257
rect -158 -325 -146 -291
rect -112 -325 -100 -291
rect -158 -359 -100 -325
rect -158 -393 -146 -359
rect -112 -393 -100 -359
rect -158 -436 -100 -393
rect 100 321 158 364
rect 100 287 112 321
rect 146 287 158 321
rect 100 253 158 287
rect 100 219 112 253
rect 146 219 158 253
rect 100 185 158 219
rect 100 151 112 185
rect 146 151 158 185
rect 100 117 158 151
rect 100 83 112 117
rect 146 83 158 117
rect 100 49 158 83
rect 100 15 112 49
rect 146 15 158 49
rect 100 -19 158 15
rect 100 -53 112 -19
rect 146 -53 158 -19
rect 100 -87 158 -53
rect 100 -121 112 -87
rect 146 -121 158 -87
rect 100 -155 158 -121
rect 100 -189 112 -155
rect 146 -189 158 -155
rect 100 -223 158 -189
rect 100 -257 112 -223
rect 146 -257 158 -223
rect 100 -291 158 -257
rect 100 -325 112 -291
rect 146 -325 158 -291
rect 100 -359 158 -325
rect 100 -393 112 -359
rect 146 -393 158 -359
rect 100 -436 158 -393
<< pdiffc >>
rect -146 287 -112 321
rect -146 219 -112 253
rect -146 151 -112 185
rect -146 83 -112 117
rect -146 15 -112 49
rect -146 -53 -112 -19
rect -146 -121 -112 -87
rect -146 -189 -112 -155
rect -146 -257 -112 -223
rect -146 -325 -112 -291
rect -146 -393 -112 -359
rect 112 287 146 321
rect 112 219 146 253
rect 112 151 146 185
rect 112 83 146 117
rect 112 15 146 49
rect 112 -53 146 -19
rect 112 -121 146 -87
rect 112 -189 146 -155
rect 112 -257 146 -223
rect 112 -325 146 -291
rect 112 -393 146 -359
<< poly >>
rect -100 445 100 461
rect -100 411 -51 445
rect -17 411 17 445
rect 51 411 100 445
rect -100 364 100 411
rect -100 -462 100 -436
<< polycont >>
rect -51 411 -17 445
rect 17 411 51 445
<< locali >>
rect -100 411 -53 445
rect -17 411 17 445
rect 53 411 100 445
rect -146 341 -112 368
rect -146 269 -112 287
rect -146 197 -112 219
rect -146 125 -112 151
rect -146 53 -112 83
rect -146 -19 -112 15
rect -146 -87 -112 -53
rect -146 -155 -112 -125
rect -146 -223 -112 -197
rect -146 -291 -112 -269
rect -146 -359 -112 -341
rect -146 -440 -112 -413
rect 112 341 146 368
rect 112 269 146 287
rect 112 197 146 219
rect 112 125 146 151
rect 112 53 146 83
rect 112 -19 146 15
rect 112 -87 146 -53
rect 112 -155 146 -125
rect 112 -223 146 -197
rect 112 -291 146 -269
rect 112 -359 146 -341
rect 112 -440 146 -413
<< viali >>
rect -53 411 -51 445
rect -51 411 -19 445
rect 19 411 51 445
rect 51 411 53 445
rect -146 321 -112 341
rect -146 307 -112 321
rect -146 253 -112 269
rect -146 235 -112 253
rect -146 185 -112 197
rect -146 163 -112 185
rect -146 117 -112 125
rect -146 91 -112 117
rect -146 49 -112 53
rect -146 19 -112 49
rect -146 -53 -112 -19
rect -146 -121 -112 -91
rect -146 -125 -112 -121
rect -146 -189 -112 -163
rect -146 -197 -112 -189
rect -146 -257 -112 -235
rect -146 -269 -112 -257
rect -146 -325 -112 -307
rect -146 -341 -112 -325
rect -146 -393 -112 -379
rect -146 -413 -112 -393
rect 112 321 146 341
rect 112 307 146 321
rect 112 253 146 269
rect 112 235 146 253
rect 112 185 146 197
rect 112 163 146 185
rect 112 117 146 125
rect 112 91 146 117
rect 112 49 146 53
rect 112 19 146 49
rect 112 -53 146 -19
rect 112 -121 146 -91
rect 112 -125 146 -121
rect 112 -189 146 -163
rect 112 -197 146 -189
rect 112 -257 146 -235
rect 112 -269 146 -257
rect 112 -325 146 -307
rect 112 -341 146 -325
rect 112 -393 146 -379
rect 112 -413 146 -393
<< metal1 >>
rect -96 445 96 451
rect -96 411 -53 445
rect -19 411 19 445
rect 53 411 96 445
rect -96 405 96 411
rect -152 341 -106 364
rect -152 307 -146 341
rect -112 307 -106 341
rect -152 269 -106 307
rect -152 235 -146 269
rect -112 235 -106 269
rect -152 197 -106 235
rect -152 163 -146 197
rect -112 163 -106 197
rect -152 125 -106 163
rect -152 91 -146 125
rect -112 91 -106 125
rect -152 53 -106 91
rect -152 19 -146 53
rect -112 19 -106 53
rect -152 -19 -106 19
rect -152 -53 -146 -19
rect -112 -53 -106 -19
rect -152 -91 -106 -53
rect -152 -125 -146 -91
rect -112 -125 -106 -91
rect -152 -163 -106 -125
rect -152 -197 -146 -163
rect -112 -197 -106 -163
rect -152 -235 -106 -197
rect -152 -269 -146 -235
rect -112 -269 -106 -235
rect -152 -307 -106 -269
rect -152 -341 -146 -307
rect -112 -341 -106 -307
rect -152 -379 -106 -341
rect -152 -413 -146 -379
rect -112 -413 -106 -379
rect -152 -436 -106 -413
rect 106 341 152 364
rect 106 307 112 341
rect 146 307 152 341
rect 106 269 152 307
rect 106 235 112 269
rect 146 235 152 269
rect 106 197 152 235
rect 106 163 112 197
rect 146 163 152 197
rect 106 125 152 163
rect 106 91 112 125
rect 146 91 152 125
rect 106 53 152 91
rect 106 19 112 53
rect 146 19 152 53
rect 106 -19 152 19
rect 106 -53 112 -19
rect 146 -53 152 -19
rect 106 -91 152 -53
rect 106 -125 112 -91
rect 146 -125 152 -91
rect 106 -163 152 -125
rect 106 -197 112 -163
rect 146 -197 152 -163
rect 106 -235 152 -197
rect 106 -269 112 -235
rect 146 -269 152 -235
rect 106 -307 152 -269
rect 106 -341 112 -307
rect 146 -341 152 -307
rect 106 -379 152 -341
rect 106 -413 112 -379
rect 146 -413 152 -379
rect 106 -436 152 -413
<< end >>
