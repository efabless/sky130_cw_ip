magic
tech sky130A
magscale 1 2
timestamp 1715625863
<< error_p >>
rect 8588 7059 11700 7121
rect 8588 6953 8650 7059
rect 8756 4446 8818 6953
rect 8756 4384 11532 4446
rect 11638 4384 11700 7059
<< nwell >>
rect 8650 6953 11638 7059
rect 8650 4384 8756 6953
rect 11532 4384 11638 6953
rect 8650 4278 11638 4384
<< nsubdiff >>
rect 8686 6989 8776 7023
rect 8810 6989 8844 7023
rect 8878 6989 8912 7023
rect 8946 6989 8980 7023
rect 9014 6989 9048 7023
rect 9082 6989 9116 7023
rect 9150 6989 9184 7023
rect 9218 6989 9252 7023
rect 9286 6989 9320 7023
rect 9354 6989 9388 7023
rect 9422 6989 9456 7023
rect 9490 6989 9524 7023
rect 9558 6989 9592 7023
rect 9626 6989 9660 7023
rect 9694 6989 9728 7023
rect 9762 6989 9796 7023
rect 9830 6989 9864 7023
rect 9898 6989 9932 7023
rect 9966 6989 10000 7023
rect 10034 6989 10068 7023
rect 10102 6989 10136 7023
rect 10170 6989 10204 7023
rect 10238 6989 10272 7023
rect 10306 6989 10340 7023
rect 10374 6989 10408 7023
rect 10442 6989 10476 7023
rect 10510 6989 10544 7023
rect 10578 6989 10612 7023
rect 10646 6989 10680 7023
rect 10714 6989 10748 7023
rect 10782 6989 10816 7023
rect 10850 6989 10884 7023
rect 10918 6989 10952 7023
rect 10986 6989 11020 7023
rect 11054 6989 11088 7023
rect 11122 6989 11156 7023
rect 11190 6989 11224 7023
rect 11258 6989 11292 7023
rect 11326 6989 11360 7023
rect 11394 6989 11428 7023
rect 11462 6989 11602 7023
rect 8686 6883 8720 6989
rect 8686 6815 8720 6849
rect 8686 6747 8720 6781
rect 8686 6679 8720 6713
rect 8686 6611 8720 6645
rect 8686 6543 8720 6577
rect 8686 6475 8720 6509
rect 8686 6407 8720 6441
rect 8686 6339 8720 6373
rect 8686 6271 8720 6305
rect 8686 6203 8720 6237
rect 8686 6135 8720 6169
rect 8686 6067 8720 6101
rect 8686 5999 8720 6033
rect 8686 5931 8720 5965
rect 8686 5863 8720 5897
rect 8686 5795 8720 5829
rect 8686 5727 8720 5761
rect 8686 5659 8720 5693
rect 8686 5591 8720 5625
rect 8686 5523 8720 5557
rect 8686 5455 8720 5489
rect 8686 5387 8720 5421
rect 8686 5319 8720 5353
rect 8686 5251 8720 5285
rect 8686 5183 8720 5217
rect 8686 5115 8720 5149
rect 8686 5047 8720 5081
rect 8686 4979 8720 5013
rect 8686 4911 8720 4945
rect 8686 4843 8720 4877
rect 8686 4775 8720 4809
rect 8686 4707 8720 4741
rect 8686 4639 8720 4673
rect 8686 4571 8720 4605
rect 8686 4503 8720 4537
rect 8686 4348 8720 4469
rect 11568 6883 11602 6989
rect 11568 6815 11602 6849
rect 11568 6747 11602 6781
rect 11568 6679 11602 6713
rect 11568 6611 11602 6645
rect 11568 6543 11602 6577
rect 11568 6475 11602 6509
rect 11568 6407 11602 6441
rect 11568 6339 11602 6373
rect 11568 6271 11602 6305
rect 11568 6203 11602 6237
rect 11568 6135 11602 6169
rect 11568 6067 11602 6101
rect 11568 5999 11602 6033
rect 11568 5931 11602 5965
rect 11568 5863 11602 5897
rect 11568 5795 11602 5829
rect 11568 5727 11602 5761
rect 11568 5659 11602 5693
rect 11568 5591 11602 5625
rect 11568 5523 11602 5557
rect 11568 5455 11602 5489
rect 11568 5387 11602 5421
rect 11568 5319 11602 5353
rect 11568 5251 11602 5285
rect 11568 5183 11602 5217
rect 11568 5115 11602 5149
rect 11568 5047 11602 5081
rect 11568 4979 11602 5013
rect 11568 4911 11602 4945
rect 11568 4843 11602 4877
rect 11568 4775 11602 4809
rect 11568 4707 11602 4741
rect 11568 4639 11602 4673
rect 11568 4571 11602 4605
rect 11568 4503 11602 4537
rect 11568 4348 11602 4469
rect 8686 4314 8844 4348
rect 8878 4314 8912 4348
rect 8946 4314 8980 4348
rect 9014 4314 9048 4348
rect 9082 4314 9116 4348
rect 9150 4314 9184 4348
rect 9218 4314 9252 4348
rect 9286 4314 9320 4348
rect 9354 4314 9388 4348
rect 9422 4314 9456 4348
rect 9490 4314 9524 4348
rect 9558 4314 9592 4348
rect 9626 4314 9660 4348
rect 9694 4314 9728 4348
rect 9762 4314 9796 4348
rect 9830 4314 9864 4348
rect 9898 4314 9932 4348
rect 9966 4314 10000 4348
rect 10034 4314 10068 4348
rect 10102 4314 10136 4348
rect 10170 4314 10204 4348
rect 10238 4314 10272 4348
rect 10306 4314 10340 4348
rect 10374 4314 10408 4348
rect 10442 4314 10476 4348
rect 10510 4314 10544 4348
rect 10578 4314 10612 4348
rect 10646 4314 10680 4348
rect 10714 4314 10748 4348
rect 10782 4314 10816 4348
rect 10850 4314 10884 4348
rect 10918 4314 10952 4348
rect 10986 4314 11020 4348
rect 11054 4314 11088 4348
rect 11122 4314 11156 4348
rect 11190 4314 11224 4348
rect 11258 4314 11292 4348
rect 11326 4314 11360 4348
rect 11394 4314 11428 4348
rect 11462 4314 11602 4348
<< nsubdiffcont >>
rect 8776 6989 8810 7023
rect 8844 6989 8878 7023
rect 8912 6989 8946 7023
rect 8980 6989 9014 7023
rect 9048 6989 9082 7023
rect 9116 6989 9150 7023
rect 9184 6989 9218 7023
rect 9252 6989 9286 7023
rect 9320 6989 9354 7023
rect 9388 6989 9422 7023
rect 9456 6989 9490 7023
rect 9524 6989 9558 7023
rect 9592 6989 9626 7023
rect 9660 6989 9694 7023
rect 9728 6989 9762 7023
rect 9796 6989 9830 7023
rect 9864 6989 9898 7023
rect 9932 6989 9966 7023
rect 10000 6989 10034 7023
rect 10068 6989 10102 7023
rect 10136 6989 10170 7023
rect 10204 6989 10238 7023
rect 10272 6989 10306 7023
rect 10340 6989 10374 7023
rect 10408 6989 10442 7023
rect 10476 6989 10510 7023
rect 10544 6989 10578 7023
rect 10612 6989 10646 7023
rect 10680 6989 10714 7023
rect 10748 6989 10782 7023
rect 10816 6989 10850 7023
rect 10884 6989 10918 7023
rect 10952 6989 10986 7023
rect 11020 6989 11054 7023
rect 11088 6989 11122 7023
rect 11156 6989 11190 7023
rect 11224 6989 11258 7023
rect 11292 6989 11326 7023
rect 11360 6989 11394 7023
rect 11428 6989 11462 7023
rect 8686 6849 8720 6883
rect 8686 6781 8720 6815
rect 8686 6713 8720 6747
rect 8686 6645 8720 6679
rect 8686 6577 8720 6611
rect 8686 6509 8720 6543
rect 8686 6441 8720 6475
rect 8686 6373 8720 6407
rect 8686 6305 8720 6339
rect 8686 6237 8720 6271
rect 8686 6169 8720 6203
rect 8686 6101 8720 6135
rect 8686 6033 8720 6067
rect 8686 5965 8720 5999
rect 8686 5897 8720 5931
rect 8686 5829 8720 5863
rect 8686 5761 8720 5795
rect 8686 5693 8720 5727
rect 8686 5625 8720 5659
rect 8686 5557 8720 5591
rect 8686 5489 8720 5523
rect 8686 5421 8720 5455
rect 8686 5353 8720 5387
rect 8686 5285 8720 5319
rect 8686 5217 8720 5251
rect 8686 5149 8720 5183
rect 8686 5081 8720 5115
rect 8686 5013 8720 5047
rect 8686 4945 8720 4979
rect 8686 4877 8720 4911
rect 8686 4809 8720 4843
rect 8686 4741 8720 4775
rect 8686 4673 8720 4707
rect 8686 4605 8720 4639
rect 8686 4537 8720 4571
rect 8686 4469 8720 4503
rect 11568 6849 11602 6883
rect 11568 6781 11602 6815
rect 11568 6713 11602 6747
rect 11568 6645 11602 6679
rect 11568 6577 11602 6611
rect 11568 6509 11602 6543
rect 11568 6441 11602 6475
rect 11568 6373 11602 6407
rect 11568 6305 11602 6339
rect 11568 6237 11602 6271
rect 11568 6169 11602 6203
rect 11568 6101 11602 6135
rect 11568 6033 11602 6067
rect 11568 5965 11602 5999
rect 11568 5897 11602 5931
rect 11568 5829 11602 5863
rect 11568 5761 11602 5795
rect 11568 5693 11602 5727
rect 11568 5625 11602 5659
rect 11568 5557 11602 5591
rect 11568 5489 11602 5523
rect 11568 5421 11602 5455
rect 11568 5353 11602 5387
rect 11568 5285 11602 5319
rect 11568 5217 11602 5251
rect 11568 5149 11602 5183
rect 11568 5081 11602 5115
rect 11568 5013 11602 5047
rect 11568 4945 11602 4979
rect 11568 4877 11602 4911
rect 11568 4809 11602 4843
rect 11568 4741 11602 4775
rect 11568 4673 11602 4707
rect 11568 4605 11602 4639
rect 11568 4537 11602 4571
rect 11568 4469 11602 4503
rect 8844 4314 8878 4348
rect 8912 4314 8946 4348
rect 8980 4314 9014 4348
rect 9048 4314 9082 4348
rect 9116 4314 9150 4348
rect 9184 4314 9218 4348
rect 9252 4314 9286 4348
rect 9320 4314 9354 4348
rect 9388 4314 9422 4348
rect 9456 4314 9490 4348
rect 9524 4314 9558 4348
rect 9592 4314 9626 4348
rect 9660 4314 9694 4348
rect 9728 4314 9762 4348
rect 9796 4314 9830 4348
rect 9864 4314 9898 4348
rect 9932 4314 9966 4348
rect 10000 4314 10034 4348
rect 10068 4314 10102 4348
rect 10136 4314 10170 4348
rect 10204 4314 10238 4348
rect 10272 4314 10306 4348
rect 10340 4314 10374 4348
rect 10408 4314 10442 4348
rect 10476 4314 10510 4348
rect 10544 4314 10578 4348
rect 10612 4314 10646 4348
rect 10680 4314 10714 4348
rect 10748 4314 10782 4348
rect 10816 4314 10850 4348
rect 10884 4314 10918 4348
rect 10952 4314 10986 4348
rect 11020 4314 11054 4348
rect 11088 4314 11122 4348
rect 11156 4314 11190 4348
rect 11224 4314 11258 4348
rect 11292 4314 11326 4348
rect 11360 4314 11394 4348
rect 11428 4314 11462 4348
<< locali >>
rect 8686 6989 8776 7023
rect 8810 6989 8844 7023
rect 8878 6989 8912 7023
rect 8946 6989 8980 7023
rect 9014 6989 9048 7023
rect 9082 6989 9116 7023
rect 9150 6989 9184 7023
rect 9218 6989 9252 7023
rect 9286 6989 9320 7023
rect 9354 6989 9388 7023
rect 9422 6989 9456 7023
rect 9490 6989 9524 7023
rect 9558 6989 9592 7023
rect 9626 6989 9660 7023
rect 9694 6989 9728 7023
rect 9762 6989 9796 7023
rect 9830 6989 9864 7023
rect 9898 6989 9932 7023
rect 9966 6989 10000 7023
rect 10034 6989 10068 7023
rect 10102 6989 10136 7023
rect 10170 6989 10204 7023
rect 10238 6989 10272 7023
rect 10306 6989 10340 7023
rect 10374 6989 10408 7023
rect 10442 6989 10476 7023
rect 10510 6989 10544 7023
rect 10578 6989 10612 7023
rect 10646 6989 10680 7023
rect 10714 6989 10748 7023
rect 10782 6989 10816 7023
rect 10850 6989 10884 7023
rect 10918 6989 10952 7023
rect 10986 6989 11020 7023
rect 11054 6989 11088 7023
rect 11122 6989 11156 7023
rect 11190 6989 11224 7023
rect 11258 6989 11292 7023
rect 11326 6989 11360 7023
rect 11394 6989 11428 7023
rect 11462 6989 11602 7023
rect 8686 6883 8720 6989
rect 8686 6815 8720 6849
rect 8686 6747 8720 6781
rect 8686 6679 8720 6713
rect 8686 6611 8720 6645
rect 8686 6543 8720 6577
rect 8686 6475 8720 6509
rect 8686 6407 8720 6441
rect 8686 6339 8720 6373
rect 8686 6271 8720 6305
rect 8686 6203 8720 6237
rect 8686 6135 8720 6169
rect 8686 6067 8720 6101
rect 8686 5999 8720 6033
rect 8686 5931 8720 5965
rect 8686 5863 8720 5897
rect 8686 5795 8720 5829
rect 8686 5727 8720 5761
rect 8686 5659 8720 5693
rect 8686 5591 8720 5625
rect 8686 5523 8720 5557
rect 8686 5455 8720 5489
rect 8686 5387 8720 5421
rect 8686 5319 8720 5353
rect 8686 5251 8720 5285
rect 8686 5183 8720 5217
rect 8686 5115 8720 5149
rect 8686 5047 8720 5081
rect 8686 4979 8720 5013
rect 8686 4911 8720 4945
rect 8686 4843 8720 4877
rect 8686 4775 8720 4809
rect 8686 4707 8720 4741
rect 8686 4639 8720 4673
rect 8686 4571 8720 4605
rect 8686 4503 8720 4537
rect 8686 4348 8720 4469
rect 11568 6883 11602 6989
rect 11568 6815 11602 6849
rect 11568 6747 11602 6781
rect 11568 6679 11602 6713
rect 11568 6611 11602 6645
rect 11568 6543 11602 6577
rect 11568 6475 11602 6509
rect 11568 6407 11602 6441
rect 11568 6339 11602 6373
rect 11568 6271 11602 6305
rect 11568 6203 11602 6237
rect 11568 6135 11602 6169
rect 11568 6067 11602 6101
rect 11568 5999 11602 6033
rect 11568 5931 11602 5965
rect 11568 5863 11602 5897
rect 11568 5795 11602 5829
rect 11568 5727 11602 5761
rect 11568 5659 11602 5693
rect 11568 5591 11602 5625
rect 11568 5523 11602 5557
rect 11568 5455 11602 5489
rect 11568 5387 11602 5421
rect 11568 5319 11602 5353
rect 11568 5251 11602 5285
rect 11568 5183 11602 5217
rect 11568 5115 11602 5149
rect 11568 5047 11602 5081
rect 11568 4979 11602 5013
rect 11568 4911 11602 4945
rect 11568 4843 11602 4877
rect 11568 4775 11602 4809
rect 11568 4707 11602 4741
rect 11568 4639 11602 4673
rect 11568 4571 11602 4605
rect 11568 4503 11602 4537
rect 11568 4348 11602 4469
rect 8686 4314 8844 4348
rect 8878 4314 8912 4348
rect 8946 4314 8980 4348
rect 9014 4314 9048 4348
rect 9082 4314 9116 4348
rect 9150 4314 9184 4348
rect 9218 4314 9252 4348
rect 9286 4314 9320 4348
rect 9354 4314 9388 4348
rect 9422 4314 9456 4348
rect 9490 4314 9524 4348
rect 9558 4314 9592 4348
rect 9626 4314 9660 4348
rect 9694 4314 9728 4348
rect 9762 4314 9796 4348
rect 9830 4314 9864 4348
rect 9898 4314 9932 4348
rect 9966 4314 10000 4348
rect 10034 4314 10068 4348
rect 10102 4314 10136 4348
rect 10170 4314 10204 4348
rect 10238 4314 10272 4348
rect 10306 4314 10340 4348
rect 10374 4314 10408 4348
rect 10442 4314 10476 4348
rect 10510 4314 10544 4348
rect 10578 4314 10612 4348
rect 10646 4314 10680 4348
rect 10714 4314 10748 4348
rect 10782 4314 10816 4348
rect 10850 4314 10884 4348
rect 10918 4314 10952 4348
rect 10986 4314 11020 4348
rect 11054 4314 11088 4348
rect 11122 4314 11156 4348
rect 11190 4314 11224 4348
rect 11258 4314 11292 4348
rect 11326 4314 11360 4348
rect 11394 4314 11428 4348
rect 11462 4314 11602 4348
<< properties >>
string path 43.250 35.030 57.925 35.030 57.925 21.655 43.515 21.655 43.515 35.030 
<< end >>
