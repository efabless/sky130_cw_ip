magic
tech sky130A
magscale 1 2
timestamp 1715010268
<< nwell >>
rect -494 -298 494 264
<< pmoslvt >>
rect -400 -236 400 164
<< pdiff >>
rect -458 151 -400 164
rect -458 117 -446 151
rect -412 117 -400 151
rect -458 83 -400 117
rect -458 49 -446 83
rect -412 49 -400 83
rect -458 15 -400 49
rect -458 -19 -446 15
rect -412 -19 -400 15
rect -458 -53 -400 -19
rect -458 -87 -446 -53
rect -412 -87 -400 -53
rect -458 -121 -400 -87
rect -458 -155 -446 -121
rect -412 -155 -400 -121
rect -458 -189 -400 -155
rect -458 -223 -446 -189
rect -412 -223 -400 -189
rect -458 -236 -400 -223
rect 400 151 458 164
rect 400 117 412 151
rect 446 117 458 151
rect 400 83 458 117
rect 400 49 412 83
rect 446 49 458 83
rect 400 15 458 49
rect 400 -19 412 15
rect 446 -19 458 15
rect 400 -53 458 -19
rect 400 -87 412 -53
rect 446 -87 458 -53
rect 400 -121 458 -87
rect 400 -155 412 -121
rect 446 -155 458 -121
rect 400 -189 458 -155
rect 400 -223 412 -189
rect 446 -223 458 -189
rect 400 -236 458 -223
<< pdiffc >>
rect -446 117 -412 151
rect -446 49 -412 83
rect -446 -19 -412 15
rect -446 -87 -412 -53
rect -446 -155 -412 -121
rect -446 -223 -412 -189
rect 412 117 446 151
rect 412 49 446 83
rect 412 -19 446 15
rect 412 -87 446 -53
rect 412 -155 446 -121
rect 412 -223 446 -189
<< poly >>
rect -400 245 400 261
rect -400 211 -357 245
rect -323 211 -289 245
rect -255 211 -221 245
rect -187 211 -153 245
rect -119 211 -85 245
rect -51 211 -17 245
rect 17 211 51 245
rect 85 211 119 245
rect 153 211 187 245
rect 221 211 255 245
rect 289 211 323 245
rect 357 211 400 245
rect -400 164 400 211
rect -400 -262 400 -236
<< polycont >>
rect -357 211 -323 245
rect -289 211 -255 245
rect -221 211 -187 245
rect -153 211 -119 245
rect -85 211 -51 245
rect -17 211 17 245
rect 51 211 85 245
rect 119 211 153 245
rect 187 211 221 245
rect 255 211 289 245
rect 323 211 357 245
<< locali >>
rect -400 211 -377 245
rect -323 211 -305 245
rect -255 211 -233 245
rect -187 211 -161 245
rect -119 211 -89 245
rect -51 211 -17 245
rect 17 211 51 245
rect 89 211 119 245
rect 161 211 187 245
rect 233 211 255 245
rect 305 211 323 245
rect 377 211 400 245
rect -446 151 -412 168
rect -446 83 -412 91
rect -446 15 -412 19
rect -446 -91 -412 -87
rect -446 -163 -412 -155
rect -446 -240 -412 -223
rect 412 151 446 168
rect 412 83 446 91
rect 412 15 446 19
rect 412 -91 446 -87
rect 412 -163 446 -155
rect 412 -240 446 -223
<< viali >>
rect -377 211 -357 245
rect -357 211 -343 245
rect -305 211 -289 245
rect -289 211 -271 245
rect -233 211 -221 245
rect -221 211 -199 245
rect -161 211 -153 245
rect -153 211 -127 245
rect -89 211 -85 245
rect -85 211 -55 245
rect -17 211 17 245
rect 55 211 85 245
rect 85 211 89 245
rect 127 211 153 245
rect 153 211 161 245
rect 199 211 221 245
rect 221 211 233 245
rect 271 211 289 245
rect 289 211 305 245
rect 343 211 357 245
rect 357 211 377 245
rect -446 117 -412 125
rect -446 91 -412 117
rect -446 49 -412 53
rect -446 19 -412 49
rect -446 -53 -412 -19
rect -446 -121 -412 -91
rect -446 -125 -412 -121
rect -446 -189 -412 -163
rect -446 -197 -412 -189
rect 412 117 446 125
rect 412 91 446 117
rect 412 49 446 53
rect 412 19 446 49
rect 412 -53 446 -19
rect 412 -121 446 -91
rect 412 -125 446 -121
rect 412 -189 446 -163
rect 412 -197 446 -189
<< metal1 >>
rect -396 245 396 251
rect -396 211 -377 245
rect -343 211 -305 245
rect -271 211 -233 245
rect -199 211 -161 245
rect -127 211 -89 245
rect -55 211 -17 245
rect 17 211 55 245
rect 89 211 127 245
rect 161 211 199 245
rect 233 211 271 245
rect 305 211 343 245
rect 377 211 396 245
rect -396 205 396 211
rect -452 125 -406 164
rect -452 91 -446 125
rect -412 91 -406 125
rect -452 53 -406 91
rect -452 19 -446 53
rect -412 19 -406 53
rect -452 -19 -406 19
rect -452 -53 -446 -19
rect -412 -53 -406 -19
rect -452 -91 -406 -53
rect -452 -125 -446 -91
rect -412 -125 -406 -91
rect -452 -163 -406 -125
rect -452 -197 -446 -163
rect -412 -197 -406 -163
rect -452 -236 -406 -197
rect 406 125 452 164
rect 406 91 412 125
rect 446 91 452 125
rect 406 53 452 91
rect 406 19 412 53
rect 446 19 452 53
rect 406 -19 452 19
rect 406 -53 412 -19
rect 446 -53 452 -19
rect 406 -91 452 -53
rect 406 -125 412 -91
rect 446 -125 452 -91
rect 406 -163 452 -125
rect 406 -197 412 -163
rect 446 -197 452 -163
rect 406 -236 452 -197
<< end >>
