magic
tech sky130A
magscale 1 2
timestamp 1715625863
<< pwell >>
rect -4272 782 4272 868
rect -4272 -782 -4186 782
rect 4186 -782 4272 782
rect -4272 -868 4272 -782
<< psubdiff >>
rect -4246 808 -4131 842
rect -4097 808 -4063 842
rect -4029 808 -3995 842
rect -3961 808 -3927 842
rect -3893 808 -3859 842
rect -3825 808 -3791 842
rect -3757 808 -3723 842
rect -3689 808 -3655 842
rect -3621 808 -3587 842
rect -3553 808 -3519 842
rect -3485 808 -3451 842
rect -3417 808 -3383 842
rect -3349 808 -3315 842
rect -3281 808 -3247 842
rect -3213 808 -3179 842
rect -3145 808 -3111 842
rect -3077 808 -3043 842
rect -3009 808 -2975 842
rect -2941 808 -2907 842
rect -2873 808 -2839 842
rect -2805 808 -2771 842
rect -2737 808 -2703 842
rect -2669 808 -2635 842
rect -2601 808 -2567 842
rect -2533 808 -2499 842
rect -2465 808 -2431 842
rect -2397 808 -2363 842
rect -2329 808 -2295 842
rect -2261 808 -2227 842
rect -2193 808 -2159 842
rect -2125 808 -2091 842
rect -2057 808 -2023 842
rect -1989 808 -1955 842
rect -1921 808 -1887 842
rect -1853 808 -1819 842
rect -1785 808 -1751 842
rect -1717 808 -1683 842
rect -1649 808 -1615 842
rect -1581 808 -1547 842
rect -1513 808 -1479 842
rect -1445 808 -1411 842
rect -1377 808 -1343 842
rect -1309 808 -1275 842
rect -1241 808 -1207 842
rect -1173 808 -1139 842
rect -1105 808 -1071 842
rect -1037 808 -1003 842
rect -969 808 -935 842
rect -901 808 -867 842
rect -833 808 -799 842
rect -765 808 -731 842
rect -697 808 -663 842
rect -629 808 -595 842
rect -561 808 -527 842
rect -493 808 -459 842
rect -425 808 -391 842
rect -357 808 -323 842
rect -289 808 -255 842
rect -221 808 -187 842
rect -153 808 -119 842
rect -85 808 -51 842
rect -17 808 17 842
rect 51 808 85 842
rect 119 808 153 842
rect 187 808 221 842
rect 255 808 289 842
rect 323 808 357 842
rect 391 808 425 842
rect 459 808 493 842
rect 527 808 561 842
rect 595 808 629 842
rect 663 808 697 842
rect 731 808 765 842
rect 799 808 833 842
rect 867 808 901 842
rect 935 808 969 842
rect 1003 808 1037 842
rect 1071 808 1105 842
rect 1139 808 1173 842
rect 1207 808 1241 842
rect 1275 808 1309 842
rect 1343 808 1377 842
rect 1411 808 1445 842
rect 1479 808 1513 842
rect 1547 808 1581 842
rect 1615 808 1649 842
rect 1683 808 1717 842
rect 1751 808 1785 842
rect 1819 808 1853 842
rect 1887 808 1921 842
rect 1955 808 1989 842
rect 2023 808 2057 842
rect 2091 808 2125 842
rect 2159 808 2193 842
rect 2227 808 2261 842
rect 2295 808 2329 842
rect 2363 808 2397 842
rect 2431 808 2465 842
rect 2499 808 2533 842
rect 2567 808 2601 842
rect 2635 808 2669 842
rect 2703 808 2737 842
rect 2771 808 2805 842
rect 2839 808 2873 842
rect 2907 808 2941 842
rect 2975 808 3009 842
rect 3043 808 3077 842
rect 3111 808 3145 842
rect 3179 808 3213 842
rect 3247 808 3281 842
rect 3315 808 3349 842
rect 3383 808 3417 842
rect 3451 808 3485 842
rect 3519 808 3553 842
rect 3587 808 3621 842
rect 3655 808 3689 842
rect 3723 808 3757 842
rect 3791 808 3825 842
rect 3859 808 3893 842
rect 3927 808 3961 842
rect 3995 808 4029 842
rect 4063 808 4097 842
rect 4131 808 4246 842
rect -4246 731 -4212 808
rect 4212 731 4246 808
rect -4246 663 -4212 697
rect -4246 595 -4212 629
rect -4246 527 -4212 561
rect -4246 459 -4212 493
rect -4246 391 -4212 425
rect -4246 323 -4212 357
rect -4246 255 -4212 289
rect -4246 187 -4212 221
rect -4246 119 -4212 153
rect -4246 51 -4212 85
rect -4246 -17 -4212 17
rect -4246 -85 -4212 -51
rect -4246 -153 -4212 -119
rect -4246 -221 -4212 -187
rect -4246 -289 -4212 -255
rect -4246 -357 -4212 -323
rect -4246 -425 -4212 -391
rect -4246 -493 -4212 -459
rect -4246 -561 -4212 -527
rect -4246 -629 -4212 -595
rect -4246 -697 -4212 -663
rect 4212 663 4246 697
rect 4212 595 4246 629
rect 4212 527 4246 561
rect 4212 459 4246 493
rect 4212 391 4246 425
rect 4212 323 4246 357
rect 4212 255 4246 289
rect 4212 187 4246 221
rect 4212 119 4246 153
rect 4212 51 4246 85
rect 4212 -17 4246 17
rect 4212 -85 4246 -51
rect 4212 -153 4246 -119
rect 4212 -221 4246 -187
rect 4212 -289 4246 -255
rect 4212 -357 4246 -323
rect 4212 -425 4246 -391
rect 4212 -493 4246 -459
rect 4212 -561 4246 -527
rect 4212 -629 4246 -595
rect 4212 -697 4246 -663
rect -4246 -808 -4212 -731
rect 4212 -808 4246 -731
rect -4246 -842 -4131 -808
rect -4097 -842 -4063 -808
rect -4029 -842 -3995 -808
rect -3961 -842 -3927 -808
rect -3893 -842 -3859 -808
rect -3825 -842 -3791 -808
rect -3757 -842 -3723 -808
rect -3689 -842 -3655 -808
rect -3621 -842 -3587 -808
rect -3553 -842 -3519 -808
rect -3485 -842 -3451 -808
rect -3417 -842 -3383 -808
rect -3349 -842 -3315 -808
rect -3281 -842 -3247 -808
rect -3213 -842 -3179 -808
rect -3145 -842 -3111 -808
rect -3077 -842 -3043 -808
rect -3009 -842 -2975 -808
rect -2941 -842 -2907 -808
rect -2873 -842 -2839 -808
rect -2805 -842 -2771 -808
rect -2737 -842 -2703 -808
rect -2669 -842 -2635 -808
rect -2601 -842 -2567 -808
rect -2533 -842 -2499 -808
rect -2465 -842 -2431 -808
rect -2397 -842 -2363 -808
rect -2329 -842 -2295 -808
rect -2261 -842 -2227 -808
rect -2193 -842 -2159 -808
rect -2125 -842 -2091 -808
rect -2057 -842 -2023 -808
rect -1989 -842 -1955 -808
rect -1921 -842 -1887 -808
rect -1853 -842 -1819 -808
rect -1785 -842 -1751 -808
rect -1717 -842 -1683 -808
rect -1649 -842 -1615 -808
rect -1581 -842 -1547 -808
rect -1513 -842 -1479 -808
rect -1445 -842 -1411 -808
rect -1377 -842 -1343 -808
rect -1309 -842 -1275 -808
rect -1241 -842 -1207 -808
rect -1173 -842 -1139 -808
rect -1105 -842 -1071 -808
rect -1037 -842 -1003 -808
rect -969 -842 -935 -808
rect -901 -842 -867 -808
rect -833 -842 -799 -808
rect -765 -842 -731 -808
rect -697 -842 -663 -808
rect -629 -842 -595 -808
rect -561 -842 -527 -808
rect -493 -842 -459 -808
rect -425 -842 -391 -808
rect -357 -842 -323 -808
rect -289 -842 -255 -808
rect -221 -842 -187 -808
rect -153 -842 -119 -808
rect -85 -842 -51 -808
rect -17 -842 17 -808
rect 51 -842 85 -808
rect 119 -842 153 -808
rect 187 -842 221 -808
rect 255 -842 289 -808
rect 323 -842 357 -808
rect 391 -842 425 -808
rect 459 -842 493 -808
rect 527 -842 561 -808
rect 595 -842 629 -808
rect 663 -842 697 -808
rect 731 -842 765 -808
rect 799 -842 833 -808
rect 867 -842 901 -808
rect 935 -842 969 -808
rect 1003 -842 1037 -808
rect 1071 -842 1105 -808
rect 1139 -842 1173 -808
rect 1207 -842 1241 -808
rect 1275 -842 1309 -808
rect 1343 -842 1377 -808
rect 1411 -842 1445 -808
rect 1479 -842 1513 -808
rect 1547 -842 1581 -808
rect 1615 -842 1649 -808
rect 1683 -842 1717 -808
rect 1751 -842 1785 -808
rect 1819 -842 1853 -808
rect 1887 -842 1921 -808
rect 1955 -842 1989 -808
rect 2023 -842 2057 -808
rect 2091 -842 2125 -808
rect 2159 -842 2193 -808
rect 2227 -842 2261 -808
rect 2295 -842 2329 -808
rect 2363 -842 2397 -808
rect 2431 -842 2465 -808
rect 2499 -842 2533 -808
rect 2567 -842 2601 -808
rect 2635 -842 2669 -808
rect 2703 -842 2737 -808
rect 2771 -842 2805 -808
rect 2839 -842 2873 -808
rect 2907 -842 2941 -808
rect 2975 -842 3009 -808
rect 3043 -842 3077 -808
rect 3111 -842 3145 -808
rect 3179 -842 3213 -808
rect 3247 -842 3281 -808
rect 3315 -842 3349 -808
rect 3383 -842 3417 -808
rect 3451 -842 3485 -808
rect 3519 -842 3553 -808
rect 3587 -842 3621 -808
rect 3655 -842 3689 -808
rect 3723 -842 3757 -808
rect 3791 -842 3825 -808
rect 3859 -842 3893 -808
rect 3927 -842 3961 -808
rect 3995 -842 4029 -808
rect 4063 -842 4097 -808
rect 4131 -842 4246 -808
<< psubdiffcont >>
rect -4131 808 -4097 842
rect -4063 808 -4029 842
rect -3995 808 -3961 842
rect -3927 808 -3893 842
rect -3859 808 -3825 842
rect -3791 808 -3757 842
rect -3723 808 -3689 842
rect -3655 808 -3621 842
rect -3587 808 -3553 842
rect -3519 808 -3485 842
rect -3451 808 -3417 842
rect -3383 808 -3349 842
rect -3315 808 -3281 842
rect -3247 808 -3213 842
rect -3179 808 -3145 842
rect -3111 808 -3077 842
rect -3043 808 -3009 842
rect -2975 808 -2941 842
rect -2907 808 -2873 842
rect -2839 808 -2805 842
rect -2771 808 -2737 842
rect -2703 808 -2669 842
rect -2635 808 -2601 842
rect -2567 808 -2533 842
rect -2499 808 -2465 842
rect -2431 808 -2397 842
rect -2363 808 -2329 842
rect -2295 808 -2261 842
rect -2227 808 -2193 842
rect -2159 808 -2125 842
rect -2091 808 -2057 842
rect -2023 808 -1989 842
rect -1955 808 -1921 842
rect -1887 808 -1853 842
rect -1819 808 -1785 842
rect -1751 808 -1717 842
rect -1683 808 -1649 842
rect -1615 808 -1581 842
rect -1547 808 -1513 842
rect -1479 808 -1445 842
rect -1411 808 -1377 842
rect -1343 808 -1309 842
rect -1275 808 -1241 842
rect -1207 808 -1173 842
rect -1139 808 -1105 842
rect -1071 808 -1037 842
rect -1003 808 -969 842
rect -935 808 -901 842
rect -867 808 -833 842
rect -799 808 -765 842
rect -731 808 -697 842
rect -663 808 -629 842
rect -595 808 -561 842
rect -527 808 -493 842
rect -459 808 -425 842
rect -391 808 -357 842
rect -323 808 -289 842
rect -255 808 -221 842
rect -187 808 -153 842
rect -119 808 -85 842
rect -51 808 -17 842
rect 17 808 51 842
rect 85 808 119 842
rect 153 808 187 842
rect 221 808 255 842
rect 289 808 323 842
rect 357 808 391 842
rect 425 808 459 842
rect 493 808 527 842
rect 561 808 595 842
rect 629 808 663 842
rect 697 808 731 842
rect 765 808 799 842
rect 833 808 867 842
rect 901 808 935 842
rect 969 808 1003 842
rect 1037 808 1071 842
rect 1105 808 1139 842
rect 1173 808 1207 842
rect 1241 808 1275 842
rect 1309 808 1343 842
rect 1377 808 1411 842
rect 1445 808 1479 842
rect 1513 808 1547 842
rect 1581 808 1615 842
rect 1649 808 1683 842
rect 1717 808 1751 842
rect 1785 808 1819 842
rect 1853 808 1887 842
rect 1921 808 1955 842
rect 1989 808 2023 842
rect 2057 808 2091 842
rect 2125 808 2159 842
rect 2193 808 2227 842
rect 2261 808 2295 842
rect 2329 808 2363 842
rect 2397 808 2431 842
rect 2465 808 2499 842
rect 2533 808 2567 842
rect 2601 808 2635 842
rect 2669 808 2703 842
rect 2737 808 2771 842
rect 2805 808 2839 842
rect 2873 808 2907 842
rect 2941 808 2975 842
rect 3009 808 3043 842
rect 3077 808 3111 842
rect 3145 808 3179 842
rect 3213 808 3247 842
rect 3281 808 3315 842
rect 3349 808 3383 842
rect 3417 808 3451 842
rect 3485 808 3519 842
rect 3553 808 3587 842
rect 3621 808 3655 842
rect 3689 808 3723 842
rect 3757 808 3791 842
rect 3825 808 3859 842
rect 3893 808 3927 842
rect 3961 808 3995 842
rect 4029 808 4063 842
rect 4097 808 4131 842
rect -4246 697 -4212 731
rect -4246 629 -4212 663
rect -4246 561 -4212 595
rect -4246 493 -4212 527
rect -4246 425 -4212 459
rect -4246 357 -4212 391
rect -4246 289 -4212 323
rect -4246 221 -4212 255
rect -4246 153 -4212 187
rect -4246 85 -4212 119
rect -4246 17 -4212 51
rect -4246 -51 -4212 -17
rect -4246 -119 -4212 -85
rect -4246 -187 -4212 -153
rect -4246 -255 -4212 -221
rect -4246 -323 -4212 -289
rect -4246 -391 -4212 -357
rect -4246 -459 -4212 -425
rect -4246 -527 -4212 -493
rect -4246 -595 -4212 -561
rect -4246 -663 -4212 -629
rect -4246 -731 -4212 -697
rect 4212 697 4246 731
rect 4212 629 4246 663
rect 4212 561 4246 595
rect 4212 493 4246 527
rect 4212 425 4246 459
rect 4212 357 4246 391
rect 4212 289 4246 323
rect 4212 221 4246 255
rect 4212 153 4246 187
rect 4212 85 4246 119
rect 4212 17 4246 51
rect 4212 -51 4246 -17
rect 4212 -119 4246 -85
rect 4212 -187 4246 -153
rect 4212 -255 4246 -221
rect 4212 -323 4246 -289
rect 4212 -391 4246 -357
rect 4212 -459 4246 -425
rect 4212 -527 4246 -493
rect 4212 -595 4246 -561
rect 4212 -663 4246 -629
rect 4212 -731 4246 -697
rect -4131 -842 -4097 -808
rect -4063 -842 -4029 -808
rect -3995 -842 -3961 -808
rect -3927 -842 -3893 -808
rect -3859 -842 -3825 -808
rect -3791 -842 -3757 -808
rect -3723 -842 -3689 -808
rect -3655 -842 -3621 -808
rect -3587 -842 -3553 -808
rect -3519 -842 -3485 -808
rect -3451 -842 -3417 -808
rect -3383 -842 -3349 -808
rect -3315 -842 -3281 -808
rect -3247 -842 -3213 -808
rect -3179 -842 -3145 -808
rect -3111 -842 -3077 -808
rect -3043 -842 -3009 -808
rect -2975 -842 -2941 -808
rect -2907 -842 -2873 -808
rect -2839 -842 -2805 -808
rect -2771 -842 -2737 -808
rect -2703 -842 -2669 -808
rect -2635 -842 -2601 -808
rect -2567 -842 -2533 -808
rect -2499 -842 -2465 -808
rect -2431 -842 -2397 -808
rect -2363 -842 -2329 -808
rect -2295 -842 -2261 -808
rect -2227 -842 -2193 -808
rect -2159 -842 -2125 -808
rect -2091 -842 -2057 -808
rect -2023 -842 -1989 -808
rect -1955 -842 -1921 -808
rect -1887 -842 -1853 -808
rect -1819 -842 -1785 -808
rect -1751 -842 -1717 -808
rect -1683 -842 -1649 -808
rect -1615 -842 -1581 -808
rect -1547 -842 -1513 -808
rect -1479 -842 -1445 -808
rect -1411 -842 -1377 -808
rect -1343 -842 -1309 -808
rect -1275 -842 -1241 -808
rect -1207 -842 -1173 -808
rect -1139 -842 -1105 -808
rect -1071 -842 -1037 -808
rect -1003 -842 -969 -808
rect -935 -842 -901 -808
rect -867 -842 -833 -808
rect -799 -842 -765 -808
rect -731 -842 -697 -808
rect -663 -842 -629 -808
rect -595 -842 -561 -808
rect -527 -842 -493 -808
rect -459 -842 -425 -808
rect -391 -842 -357 -808
rect -323 -842 -289 -808
rect -255 -842 -221 -808
rect -187 -842 -153 -808
rect -119 -842 -85 -808
rect -51 -842 -17 -808
rect 17 -842 51 -808
rect 85 -842 119 -808
rect 153 -842 187 -808
rect 221 -842 255 -808
rect 289 -842 323 -808
rect 357 -842 391 -808
rect 425 -842 459 -808
rect 493 -842 527 -808
rect 561 -842 595 -808
rect 629 -842 663 -808
rect 697 -842 731 -808
rect 765 -842 799 -808
rect 833 -842 867 -808
rect 901 -842 935 -808
rect 969 -842 1003 -808
rect 1037 -842 1071 -808
rect 1105 -842 1139 -808
rect 1173 -842 1207 -808
rect 1241 -842 1275 -808
rect 1309 -842 1343 -808
rect 1377 -842 1411 -808
rect 1445 -842 1479 -808
rect 1513 -842 1547 -808
rect 1581 -842 1615 -808
rect 1649 -842 1683 -808
rect 1717 -842 1751 -808
rect 1785 -842 1819 -808
rect 1853 -842 1887 -808
rect 1921 -842 1955 -808
rect 1989 -842 2023 -808
rect 2057 -842 2091 -808
rect 2125 -842 2159 -808
rect 2193 -842 2227 -808
rect 2261 -842 2295 -808
rect 2329 -842 2363 -808
rect 2397 -842 2431 -808
rect 2465 -842 2499 -808
rect 2533 -842 2567 -808
rect 2601 -842 2635 -808
rect 2669 -842 2703 -808
rect 2737 -842 2771 -808
rect 2805 -842 2839 -808
rect 2873 -842 2907 -808
rect 2941 -842 2975 -808
rect 3009 -842 3043 -808
rect 3077 -842 3111 -808
rect 3145 -842 3179 -808
rect 3213 -842 3247 -808
rect 3281 -842 3315 -808
rect 3349 -842 3383 -808
rect 3417 -842 3451 -808
rect 3485 -842 3519 -808
rect 3553 -842 3587 -808
rect 3621 -842 3655 -808
rect 3689 -842 3723 -808
rect 3757 -842 3791 -808
rect 3825 -842 3859 -808
rect 3893 -842 3927 -808
rect 3961 -842 3995 -808
rect 4029 -842 4063 -808
rect 4097 -842 4131 -808
<< xpolycontact >>
rect -4116 276 -3834 712
rect -4116 -712 -3834 -276
rect -3586 276 -3304 712
rect -3586 -712 -3304 -276
rect -3056 276 -2774 712
rect -3056 -712 -2774 -276
rect -2526 276 -2244 712
rect -2526 -712 -2244 -276
rect -1996 276 -1714 712
rect -1996 -712 -1714 -276
rect -1466 276 -1184 712
rect -1466 -712 -1184 -276
rect -936 276 -654 712
rect -936 -712 -654 -276
rect -406 276 -124 712
rect -406 -712 -124 -276
rect 124 276 406 712
rect 124 -712 406 -276
rect 654 276 936 712
rect 654 -712 936 -276
rect 1184 276 1466 712
rect 1184 -712 1466 -276
rect 1714 276 1996 712
rect 1714 -712 1996 -276
rect 2244 276 2526 712
rect 2244 -712 2526 -276
rect 2774 276 3056 712
rect 2774 -712 3056 -276
rect 3304 276 3586 712
rect 3304 -712 3586 -276
rect 3834 276 4116 712
rect 3834 -712 4116 -276
<< ppolyres >>
rect -4116 -276 -3834 276
rect -3586 -276 -3304 276
rect -3056 -276 -2774 276
rect -2526 -276 -2244 276
rect -1996 -276 -1714 276
rect -1466 -276 -1184 276
rect -936 -276 -654 276
rect -406 -276 -124 276
rect 124 -276 406 276
rect 654 -276 936 276
rect 1184 -276 1466 276
rect 1714 -276 1996 276
rect 2244 -276 2526 276
rect 2774 -276 3056 276
rect 3304 -276 3586 276
rect 3834 -276 4116 276
<< locali >>
rect -4246 808 -4131 842
rect -4097 808 -4063 842
rect -4029 808 -3995 842
rect -3961 808 -3927 842
rect -3893 808 -3859 842
rect -3825 808 -3791 842
rect -3757 808 -3723 842
rect -3689 808 -3655 842
rect -3621 808 -3587 842
rect -3553 808 -3519 842
rect -3485 808 -3451 842
rect -3417 808 -3383 842
rect -3349 808 -3315 842
rect -3281 808 -3247 842
rect -3213 808 -3179 842
rect -3145 808 -3111 842
rect -3077 808 -3043 842
rect -3009 808 -2975 842
rect -2941 808 -2907 842
rect -2873 808 -2839 842
rect -2805 808 -2771 842
rect -2737 808 -2703 842
rect -2669 808 -2635 842
rect -2601 808 -2567 842
rect -2533 808 -2499 842
rect -2465 808 -2431 842
rect -2397 808 -2363 842
rect -2329 808 -2295 842
rect -2261 808 -2227 842
rect -2193 808 -2159 842
rect -2125 808 -2091 842
rect -2057 808 -2023 842
rect -1989 808 -1955 842
rect -1921 808 -1887 842
rect -1853 808 -1819 842
rect -1785 808 -1751 842
rect -1717 808 -1683 842
rect -1649 808 -1615 842
rect -1581 808 -1547 842
rect -1513 808 -1479 842
rect -1445 808 -1411 842
rect -1377 808 -1343 842
rect -1309 808 -1275 842
rect -1241 808 -1207 842
rect -1173 808 -1139 842
rect -1105 808 -1071 842
rect -1037 808 -1003 842
rect -969 808 -935 842
rect -901 808 -867 842
rect -833 808 -799 842
rect -765 808 -731 842
rect -697 808 -663 842
rect -629 808 -595 842
rect -561 808 -527 842
rect -493 808 -459 842
rect -425 808 -391 842
rect -357 808 -323 842
rect -289 808 -255 842
rect -221 808 -187 842
rect -153 808 -119 842
rect -85 808 -51 842
rect -17 808 17 842
rect 51 808 85 842
rect 119 808 153 842
rect 187 808 221 842
rect 255 808 289 842
rect 323 808 357 842
rect 391 808 425 842
rect 459 808 493 842
rect 527 808 561 842
rect 595 808 629 842
rect 663 808 697 842
rect 731 808 765 842
rect 799 808 833 842
rect 867 808 901 842
rect 935 808 969 842
rect 1003 808 1037 842
rect 1071 808 1105 842
rect 1139 808 1173 842
rect 1207 808 1241 842
rect 1275 808 1309 842
rect 1343 808 1377 842
rect 1411 808 1445 842
rect 1479 808 1513 842
rect 1547 808 1581 842
rect 1615 808 1649 842
rect 1683 808 1717 842
rect 1751 808 1785 842
rect 1819 808 1853 842
rect 1887 808 1921 842
rect 1955 808 1989 842
rect 2023 808 2057 842
rect 2091 808 2125 842
rect 2159 808 2193 842
rect 2227 808 2261 842
rect 2295 808 2329 842
rect 2363 808 2397 842
rect 2431 808 2465 842
rect 2499 808 2533 842
rect 2567 808 2601 842
rect 2635 808 2669 842
rect 2703 808 2737 842
rect 2771 808 2805 842
rect 2839 808 2873 842
rect 2907 808 2941 842
rect 2975 808 3009 842
rect 3043 808 3077 842
rect 3111 808 3145 842
rect 3179 808 3213 842
rect 3247 808 3281 842
rect 3315 808 3349 842
rect 3383 808 3417 842
rect 3451 808 3485 842
rect 3519 808 3553 842
rect 3587 808 3621 842
rect 3655 808 3689 842
rect 3723 808 3757 842
rect 3791 808 3825 842
rect 3859 808 3893 842
rect 3927 808 3961 842
rect 3995 808 4029 842
rect 4063 808 4097 842
rect 4131 808 4246 842
rect -4246 731 -4212 808
rect 4212 731 4246 808
rect -4246 663 -4212 697
rect -4246 595 -4212 629
rect -4246 527 -4212 561
rect -4246 459 -4212 493
rect -4246 391 -4212 425
rect -4246 323 -4212 357
rect -4246 255 -4212 289
rect 4212 663 4246 697
rect 4212 595 4246 629
rect 4212 527 4246 561
rect 4212 459 4246 493
rect 4212 391 4246 425
rect 4212 323 4246 357
rect -4246 187 -4212 221
rect -4246 119 -4212 153
rect -4246 51 -4212 85
rect -4246 -17 -4212 17
rect -4246 -85 -4212 -51
rect -4246 -153 -4212 -119
rect -4246 -221 -4212 -187
rect -4246 -289 -4212 -255
rect 4212 255 4246 289
rect 4212 187 4246 221
rect 4212 119 4246 153
rect 4212 51 4246 85
rect 4212 -17 4246 17
rect 4212 -85 4246 -51
rect 4212 -153 4246 -119
rect 4212 -221 4246 -187
rect -4246 -357 -4212 -323
rect -4246 -425 -4212 -391
rect -4246 -493 -4212 -459
rect -4246 -561 -4212 -527
rect -4246 -629 -4212 -595
rect -4246 -697 -4212 -663
rect 4212 -289 4246 -255
rect 4212 -357 4246 -323
rect 4212 -425 4246 -391
rect 4212 -493 4246 -459
rect 4212 -561 4246 -527
rect 4212 -629 4246 -595
rect 4212 -697 4246 -663
rect -4246 -808 -4212 -731
rect 4212 -808 4246 -731
rect -4246 -842 -4131 -808
rect -4097 -842 -4063 -808
rect -4029 -842 -3995 -808
rect -3961 -842 -3927 -808
rect -3893 -842 -3859 -808
rect -3825 -842 -3791 -808
rect -3757 -842 -3723 -808
rect -3689 -842 -3655 -808
rect -3621 -842 -3587 -808
rect -3553 -842 -3519 -808
rect -3485 -842 -3451 -808
rect -3417 -842 -3383 -808
rect -3349 -842 -3315 -808
rect -3281 -842 -3247 -808
rect -3213 -842 -3179 -808
rect -3145 -842 -3111 -808
rect -3077 -842 -3043 -808
rect -3009 -842 -2975 -808
rect -2941 -842 -2907 -808
rect -2873 -842 -2839 -808
rect -2805 -842 -2771 -808
rect -2737 -842 -2703 -808
rect -2669 -842 -2635 -808
rect -2601 -842 -2567 -808
rect -2533 -842 -2499 -808
rect -2465 -842 -2431 -808
rect -2397 -842 -2363 -808
rect -2329 -842 -2295 -808
rect -2261 -842 -2227 -808
rect -2193 -842 -2159 -808
rect -2125 -842 -2091 -808
rect -2057 -842 -2023 -808
rect -1989 -842 -1955 -808
rect -1921 -842 -1887 -808
rect -1853 -842 -1819 -808
rect -1785 -842 -1751 -808
rect -1717 -842 -1683 -808
rect -1649 -842 -1615 -808
rect -1581 -842 -1547 -808
rect -1513 -842 -1479 -808
rect -1445 -842 -1411 -808
rect -1377 -842 -1343 -808
rect -1309 -842 -1275 -808
rect -1241 -842 -1207 -808
rect -1173 -842 -1139 -808
rect -1105 -842 -1071 -808
rect -1037 -842 -1003 -808
rect -969 -842 -935 -808
rect -901 -842 -867 -808
rect -833 -842 -799 -808
rect -765 -842 -731 -808
rect -697 -842 -663 -808
rect -629 -842 -595 -808
rect -561 -842 -527 -808
rect -493 -842 -459 -808
rect -425 -842 -391 -808
rect -357 -842 -323 -808
rect -289 -842 -255 -808
rect -221 -842 -187 -808
rect -153 -842 -119 -808
rect -85 -842 -51 -808
rect -17 -842 17 -808
rect 51 -842 85 -808
rect 119 -842 153 -808
rect 187 -842 221 -808
rect 255 -842 289 -808
rect 323 -842 357 -808
rect 391 -842 425 -808
rect 459 -842 493 -808
rect 527 -842 561 -808
rect 595 -842 629 -808
rect 663 -842 697 -808
rect 731 -842 765 -808
rect 799 -842 833 -808
rect 867 -842 901 -808
rect 935 -842 969 -808
rect 1003 -842 1037 -808
rect 1071 -842 1105 -808
rect 1139 -842 1173 -808
rect 1207 -842 1241 -808
rect 1275 -842 1309 -808
rect 1343 -842 1377 -808
rect 1411 -842 1445 -808
rect 1479 -842 1513 -808
rect 1547 -842 1581 -808
rect 1615 -842 1649 -808
rect 1683 -842 1717 -808
rect 1751 -842 1785 -808
rect 1819 -842 1853 -808
rect 1887 -842 1921 -808
rect 1955 -842 1989 -808
rect 2023 -842 2057 -808
rect 2091 -842 2125 -808
rect 2159 -842 2193 -808
rect 2227 -842 2261 -808
rect 2295 -842 2329 -808
rect 2363 -842 2397 -808
rect 2431 -842 2465 -808
rect 2499 -842 2533 -808
rect 2567 -842 2601 -808
rect 2635 -842 2669 -808
rect 2703 -842 2737 -808
rect 2771 -842 2805 -808
rect 2839 -842 2873 -808
rect 2907 -842 2941 -808
rect 2975 -842 3009 -808
rect 3043 -842 3077 -808
rect 3111 -842 3145 -808
rect 3179 -842 3213 -808
rect 3247 -842 3281 -808
rect 3315 -842 3349 -808
rect 3383 -842 3417 -808
rect 3451 -842 3485 -808
rect 3519 -842 3553 -808
rect 3587 -842 3621 -808
rect 3655 -842 3689 -808
rect 3723 -842 3757 -808
rect 3791 -842 3825 -808
rect 3859 -842 3893 -808
rect 3927 -842 3961 -808
rect 3995 -842 4029 -808
rect 4063 -842 4097 -808
rect 4131 -842 4246 -808
<< viali >>
rect -4100 298 -3850 692
rect -3570 298 -3320 692
rect -3040 298 -2790 692
rect -2510 298 -2260 692
rect -1980 298 -1730 692
rect -1450 298 -1200 692
rect -920 298 -670 692
rect -390 298 -140 692
rect 140 298 390 692
rect 670 298 920 692
rect 1200 298 1450 692
rect 1730 298 1980 692
rect 2260 298 2510 692
rect 2790 298 3040 692
rect 3320 298 3570 692
rect 3850 298 4100 692
rect -4100 -693 -3850 -299
rect -3570 -693 -3320 -299
rect -3040 -693 -2790 -299
rect -2510 -693 -2260 -299
rect -1980 -693 -1730 -299
rect -1450 -693 -1200 -299
rect -920 -693 -670 -299
rect -390 -693 -140 -299
rect 140 -693 390 -299
rect 670 -693 920 -299
rect 1200 -693 1450 -299
rect 1730 -693 1980 -299
rect 2260 -693 2510 -299
rect 2790 -693 3040 -299
rect 3320 -693 3570 -299
rect 3850 -693 4100 -299
<< metal1 >>
rect -4106 692 -3844 706
rect -4106 298 -4100 692
rect -3850 298 -3844 692
rect -4106 285 -3844 298
rect -3576 692 -3314 706
rect -3576 298 -3570 692
rect -3320 298 -3314 692
rect -3576 285 -3314 298
rect -3046 692 -2784 706
rect -3046 298 -3040 692
rect -2790 298 -2784 692
rect -3046 285 -2784 298
rect -2516 692 -2254 706
rect -2516 298 -2510 692
rect -2260 298 -2254 692
rect -2516 285 -2254 298
rect -1986 692 -1724 706
rect -1986 298 -1980 692
rect -1730 298 -1724 692
rect -1986 285 -1724 298
rect -1456 692 -1194 706
rect -1456 298 -1450 692
rect -1200 298 -1194 692
rect -1456 285 -1194 298
rect -926 692 -664 706
rect -926 298 -920 692
rect -670 298 -664 692
rect -926 285 -664 298
rect -396 692 -134 706
rect -396 298 -390 692
rect -140 298 -134 692
rect -396 285 -134 298
rect 134 692 396 706
rect 134 298 140 692
rect 390 298 396 692
rect 134 285 396 298
rect 664 692 926 706
rect 664 298 670 692
rect 920 298 926 692
rect 664 285 926 298
rect 1194 692 1456 706
rect 1194 298 1200 692
rect 1450 298 1456 692
rect 1194 285 1456 298
rect 1724 692 1986 706
rect 1724 298 1730 692
rect 1980 298 1986 692
rect 1724 285 1986 298
rect 2254 692 2516 706
rect 2254 298 2260 692
rect 2510 298 2516 692
rect 2254 285 2516 298
rect 2784 692 3046 706
rect 2784 298 2790 692
rect 3040 298 3046 692
rect 2784 285 3046 298
rect 3314 692 3576 706
rect 3314 298 3320 692
rect 3570 298 3576 692
rect 3314 285 3576 298
rect 3844 692 4106 706
rect 3844 298 3850 692
rect 4100 298 4106 692
rect 3844 285 4106 298
rect -4106 -299 -3844 -285
rect -4106 -693 -4100 -299
rect -3850 -693 -3844 -299
rect -4106 -706 -3844 -693
rect -3576 -299 -3314 -285
rect -3576 -693 -3570 -299
rect -3320 -693 -3314 -299
rect -3576 -706 -3314 -693
rect -3046 -299 -2784 -285
rect -3046 -693 -3040 -299
rect -2790 -693 -2784 -299
rect -3046 -706 -2784 -693
rect -2516 -299 -2254 -285
rect -2516 -693 -2510 -299
rect -2260 -693 -2254 -299
rect -2516 -706 -2254 -693
rect -1986 -299 -1724 -285
rect -1986 -693 -1980 -299
rect -1730 -693 -1724 -299
rect -1986 -706 -1724 -693
rect -1456 -299 -1194 -285
rect -1456 -693 -1450 -299
rect -1200 -693 -1194 -299
rect -1456 -706 -1194 -693
rect -926 -299 -664 -285
rect -926 -693 -920 -299
rect -670 -693 -664 -299
rect -926 -706 -664 -693
rect -396 -299 -134 -285
rect -396 -693 -390 -299
rect -140 -693 -134 -299
rect -396 -706 -134 -693
rect 134 -299 396 -285
rect 134 -693 140 -299
rect 390 -693 396 -299
rect 134 -706 396 -693
rect 664 -299 926 -285
rect 664 -693 670 -299
rect 920 -693 926 -299
rect 664 -706 926 -693
rect 1194 -299 1456 -285
rect 1194 -693 1200 -299
rect 1450 -693 1456 -299
rect 1194 -706 1456 -693
rect 1724 -299 1986 -285
rect 1724 -693 1730 -299
rect 1980 -693 1986 -299
rect 1724 -706 1986 -693
rect 2254 -299 2516 -285
rect 2254 -693 2260 -299
rect 2510 -693 2516 -299
rect 2254 -706 2516 -693
rect 2784 -299 3046 -285
rect 2784 -693 2790 -299
rect 3040 -693 3046 -299
rect 2784 -706 3046 -693
rect 3314 -299 3576 -285
rect 3314 -693 3320 -299
rect 3570 -693 3576 -299
rect 3314 -706 3576 -693
rect 3844 -299 4106 -285
rect 3844 -693 3850 -299
rect 4100 -693 4106 -299
rect 3844 -706 4106 -693
<< properties >>
string FIXED_BBOX -4229 -825 4229 825
<< end >>
