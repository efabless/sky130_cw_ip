magic
tech sky130A
magscale 1 2
timestamp 1715010268
<< error_p >>
rect 60 730 94 736
rect 60 708 66 730
rect 88 708 94 730
rect 60 702 94 708
rect 132 730 166 736
rect 132 708 138 730
rect 160 708 166 730
rect 132 702 166 708
rect 204 730 238 736
rect 204 708 210 730
rect 232 708 238 730
rect 204 702 238 708
rect 276 730 310 736
rect 276 708 282 730
rect 304 708 310 730
rect 276 702 310 708
rect 486 730 520 736
rect 486 708 492 730
rect 514 708 520 730
rect 486 702 520 708
rect 558 730 592 736
rect 558 708 564 730
rect 586 708 592 730
rect 558 702 592 708
rect 630 730 664 736
rect 630 708 636 730
rect 658 708 664 730
rect 630 702 664 708
rect 702 730 736 736
rect 702 708 708 730
rect 730 708 736 730
rect 702 702 736 708
rect 60 658 94 664
rect 60 636 66 658
rect 88 636 94 658
rect 60 630 94 636
rect 702 658 736 664
rect 702 636 708 658
rect 730 636 736 658
rect 702 630 736 636
rect 60 586 94 592
rect 60 564 66 586
rect 88 564 94 586
rect 60 558 94 564
rect 208 582 242 588
rect 208 560 214 582
rect 236 560 242 582
rect 208 554 242 560
rect 280 582 314 588
rect 280 560 286 582
rect 308 560 314 582
rect 280 554 314 560
rect 482 582 516 588
rect 482 560 488 582
rect 510 560 516 582
rect 482 554 516 560
rect 554 582 588 588
rect 554 560 560 582
rect 582 560 588 582
rect 554 554 588 560
rect 702 586 736 592
rect 702 564 708 586
rect 730 564 736 586
rect 702 558 736 564
rect 60 514 94 520
rect 60 492 66 514
rect 88 492 94 514
rect 60 486 94 492
rect 208 510 242 516
rect 208 488 214 510
rect 236 488 242 510
rect 208 482 242 488
rect 554 510 588 516
rect 554 488 560 510
rect 582 488 588 510
rect 554 482 588 488
rect 702 514 736 520
rect 702 492 708 514
rect 730 492 736 514
rect 702 486 736 492
rect 60 304 94 310
rect 60 282 66 304
rect 88 282 94 304
rect 60 276 94 282
rect 208 308 242 314
rect 208 286 214 308
rect 236 286 242 308
rect 208 280 242 286
rect 554 308 588 314
rect 554 286 560 308
rect 582 286 588 308
rect 554 280 588 286
rect 702 304 736 310
rect 702 282 708 304
rect 730 282 736 304
rect 702 276 736 282
rect 60 232 94 238
rect 60 210 66 232
rect 88 210 94 232
rect 60 204 94 210
rect 208 236 242 242
rect 208 214 214 236
rect 236 214 242 236
rect 208 208 242 214
rect 280 236 314 242
rect 280 214 286 236
rect 308 214 314 236
rect 280 208 314 214
rect 482 236 516 242
rect 482 214 488 236
rect 510 214 516 236
rect 482 208 516 214
rect 554 236 588 242
rect 554 214 560 236
rect 582 214 588 236
rect 554 208 588 214
rect 702 232 736 238
rect 702 210 708 232
rect 730 210 736 232
rect 702 204 736 210
rect 60 160 94 166
rect 60 138 66 160
rect 88 138 94 160
rect 60 132 94 138
rect 702 160 736 166
rect 702 138 708 160
rect 730 138 736 160
rect 702 132 736 138
rect 60 88 94 94
rect 60 66 66 88
rect 88 66 94 88
rect 60 60 94 66
rect 132 88 166 94
rect 132 66 138 88
rect 160 66 166 88
rect 132 60 166 66
rect 204 88 238 94
rect 204 66 210 88
rect 232 66 238 88
rect 204 60 238 66
rect 276 88 310 94
rect 276 66 282 88
rect 304 66 310 88
rect 276 60 310 66
rect 486 88 520 94
rect 486 66 492 88
rect 514 66 520 88
rect 486 60 520 66
rect 558 88 592 94
rect 558 66 564 88
rect 586 66 592 88
rect 558 60 592 66
rect 630 88 664 94
rect 630 66 636 88
rect 658 66 664 88
rect 630 60 664 66
rect 702 88 736 94
rect 702 66 708 88
rect 730 66 736 88
rect 702 60 736 66
<< pwell >>
rect 0 643 796 796
rect 0 153 153 643
rect 643 153 796 643
rect 0 0 796 153
<< nbase >>
rect 153 153 643 643
<< pdiff >>
rect 330 449 466 466
rect 330 347 347 449
rect 449 347 466 449
rect 330 330 466 347
<< pdiffc >>
rect 347 347 449 449
<< psubdiff >>
rect 26 736 770 770
rect 26 702 60 736
rect 94 702 128 736
rect 162 702 196 736
rect 230 702 264 736
rect 298 702 498 736
rect 532 702 566 736
rect 600 702 634 736
rect 668 702 702 736
rect 736 702 770 736
rect 26 669 770 702
rect 26 668 127 669
rect 26 634 60 668
rect 94 634 127 668
rect 26 600 127 634
rect 669 668 770 669
rect 669 634 702 668
rect 736 634 770 668
rect 26 566 60 600
rect 94 566 127 600
rect 26 532 127 566
rect 26 498 60 532
rect 94 498 127 532
rect 26 298 127 498
rect 26 264 60 298
rect 94 264 127 298
rect 26 230 127 264
rect 26 196 60 230
rect 94 196 127 230
rect 26 162 127 196
rect 669 600 770 634
rect 669 566 702 600
rect 736 566 770 600
rect 669 532 770 566
rect 669 498 702 532
rect 736 498 770 532
rect 669 298 770 498
rect 669 264 702 298
rect 736 264 770 298
rect 669 230 770 264
rect 669 196 702 230
rect 736 196 770 230
rect 26 128 60 162
rect 94 128 127 162
rect 26 127 127 128
rect 669 162 770 196
rect 669 128 702 162
rect 736 128 770 162
rect 669 127 770 128
rect 26 94 770 127
rect 26 60 60 94
rect 94 60 128 94
rect 162 60 196 94
rect 230 60 264 94
rect 298 60 498 94
rect 532 60 566 94
rect 600 60 634 94
rect 668 60 702 94
rect 736 60 770 94
rect 26 26 770 60
<< nsubdiff >>
rect 189 583 607 607
rect 189 549 213 583
rect 247 549 281 583
rect 315 549 481 583
rect 515 549 549 583
rect 583 549 607 583
rect 189 535 607 549
rect 189 515 261 535
rect 189 481 213 515
rect 247 481 261 515
rect 189 315 261 481
rect 535 515 607 535
rect 535 481 549 515
rect 583 481 607 515
rect 189 281 213 315
rect 247 281 261 315
rect 189 261 261 281
rect 535 315 607 481
rect 535 281 549 315
rect 583 281 607 315
rect 535 261 607 281
rect 189 247 607 261
rect 189 213 213 247
rect 247 213 281 247
rect 315 213 481 247
rect 515 213 549 247
rect 583 213 607 247
rect 189 189 607 213
<< psubdiffcont >>
rect 60 702 94 736
rect 128 702 162 736
rect 196 702 230 736
rect 264 702 298 736
rect 498 702 532 736
rect 566 702 600 736
rect 634 702 668 736
rect 702 702 736 736
rect 60 634 94 668
rect 702 634 736 668
rect 60 566 94 600
rect 60 498 94 532
rect 60 264 94 298
rect 60 196 94 230
rect 702 566 736 600
rect 702 498 736 532
rect 702 264 736 298
rect 702 196 736 230
rect 60 128 94 162
rect 702 128 736 162
rect 60 60 94 94
rect 128 60 162 94
rect 196 60 230 94
rect 264 60 298 94
rect 498 60 532 94
rect 566 60 600 94
rect 634 60 668 94
rect 702 60 736 94
<< nsubdiffcont >>
rect 213 549 247 583
rect 281 549 315 583
rect 481 549 515 583
rect 549 549 583 583
rect 213 481 247 515
rect 549 481 583 515
rect 213 281 247 315
rect 549 281 583 315
rect 213 213 247 247
rect 281 213 315 247
rect 481 213 515 247
rect 549 213 583 247
<< locali >>
rect 26 736 770 770
rect 26 702 60 736
rect 94 702 128 736
rect 166 702 196 736
rect 238 702 264 736
rect 310 702 486 736
rect 532 702 558 736
rect 600 702 630 736
rect 668 702 702 736
rect 736 702 770 736
rect 26 669 770 702
rect 26 668 127 669
rect 26 630 60 668
rect 94 630 127 668
rect 26 600 127 630
rect 669 668 770 669
rect 669 630 702 668
rect 736 630 770 668
rect 26 558 60 600
rect 94 558 127 600
rect 26 532 127 558
rect 26 486 60 532
rect 94 486 127 532
rect 26 310 127 486
rect 26 264 60 310
rect 94 264 127 310
rect 26 238 127 264
rect 26 196 60 238
rect 94 196 127 238
rect 26 166 127 196
rect 189 588 607 607
rect 189 554 208 588
rect 242 583 280 588
rect 314 583 482 588
rect 516 583 554 588
rect 247 554 280 583
rect 189 549 213 554
rect 247 549 281 554
rect 315 549 481 583
rect 516 554 549 583
rect 588 554 607 588
rect 515 549 549 554
rect 583 549 607 554
rect 189 535 607 549
rect 189 516 261 535
rect 189 482 208 516
rect 242 515 261 516
rect 189 481 213 482
rect 247 481 261 515
rect 189 315 261 481
rect 535 516 607 535
rect 535 515 554 516
rect 535 481 549 515
rect 588 482 607 516
rect 583 481 607 482
rect 319 463 477 477
rect 319 429 333 463
rect 367 449 429 463
rect 463 429 477 463
rect 319 367 347 429
rect 449 367 477 429
rect 319 333 333 367
rect 367 333 429 347
rect 463 333 477 367
rect 319 319 477 333
rect 189 314 213 315
rect 189 280 208 314
rect 247 281 261 315
rect 242 280 261 281
rect 189 261 261 280
rect 535 315 607 481
rect 535 281 549 315
rect 583 314 607 315
rect 535 280 554 281
rect 588 280 607 314
rect 535 261 607 280
rect 189 247 607 261
rect 189 242 213 247
rect 247 242 281 247
rect 189 208 208 242
rect 247 213 280 242
rect 315 213 481 247
rect 515 242 549 247
rect 583 242 607 247
rect 516 213 549 242
rect 242 208 280 213
rect 314 208 482 213
rect 516 208 554 213
rect 588 208 607 242
rect 189 189 607 208
rect 669 600 770 630
rect 669 558 702 600
rect 736 558 770 600
rect 669 532 770 558
rect 669 486 702 532
rect 736 486 770 532
rect 669 310 770 486
rect 669 264 702 310
rect 736 264 770 310
rect 669 238 770 264
rect 669 196 702 238
rect 736 196 770 238
rect 26 128 60 166
rect 94 128 127 166
rect 26 127 127 128
rect 669 166 770 196
rect 669 128 702 166
rect 736 128 770 166
rect 669 127 770 128
rect 26 94 770 127
rect 26 60 60 94
rect 94 60 128 94
rect 166 60 196 94
rect 238 60 264 94
rect 310 60 486 94
rect 532 60 558 94
rect 600 60 630 94
rect 668 60 702 94
rect 736 60 770 94
rect 26 26 770 60
<< viali >>
rect 60 702 94 736
rect 132 702 162 736
rect 162 702 166 736
rect 204 702 230 736
rect 230 702 238 736
rect 276 702 298 736
rect 298 702 310 736
rect 486 702 498 736
rect 498 702 520 736
rect 558 702 566 736
rect 566 702 592 736
rect 630 702 634 736
rect 634 702 664 736
rect 702 702 736 736
rect 60 634 94 664
rect 60 630 94 634
rect 702 634 736 664
rect 702 630 736 634
rect 60 566 94 592
rect 60 558 94 566
rect 60 498 94 520
rect 60 486 94 498
rect 60 298 94 310
rect 60 276 94 298
rect 60 230 94 238
rect 60 204 94 230
rect 208 583 242 588
rect 280 583 314 588
rect 482 583 516 588
rect 554 583 588 588
rect 208 554 213 583
rect 213 554 242 583
rect 280 554 281 583
rect 281 554 314 583
rect 482 554 515 583
rect 515 554 516 583
rect 554 554 583 583
rect 583 554 588 583
rect 208 515 242 516
rect 208 482 213 515
rect 213 482 242 515
rect 554 515 588 516
rect 554 482 583 515
rect 583 482 588 515
rect 333 449 367 463
rect 429 449 463 463
rect 333 429 347 449
rect 347 429 367 449
rect 429 429 449 449
rect 449 429 463 449
rect 333 347 347 367
rect 347 347 367 367
rect 429 347 449 367
rect 449 347 463 367
rect 333 333 367 347
rect 429 333 463 347
rect 208 281 213 314
rect 213 281 242 314
rect 208 280 242 281
rect 554 281 583 314
rect 583 281 588 314
rect 554 280 588 281
rect 208 213 213 242
rect 213 213 242 242
rect 280 213 281 242
rect 281 213 314 242
rect 482 213 515 242
rect 515 213 516 242
rect 554 213 583 242
rect 583 213 588 242
rect 208 208 242 213
rect 280 208 314 213
rect 482 208 516 213
rect 554 208 588 213
rect 702 566 736 592
rect 702 558 736 566
rect 702 498 736 520
rect 702 486 736 498
rect 702 298 736 310
rect 702 276 736 298
rect 702 230 736 238
rect 702 204 736 230
rect 60 162 94 166
rect 60 132 94 162
rect 702 162 736 166
rect 702 132 736 162
rect 60 60 94 94
rect 132 60 162 94
rect 162 60 166 94
rect 204 60 230 94
rect 230 60 238 94
rect 276 60 298 94
rect 298 60 310 94
rect 486 60 498 94
rect 498 60 520 94
rect 558 60 566 94
rect 566 60 592 94
rect 630 60 634 94
rect 634 60 664 94
rect 702 60 736 94
<< metal1 >>
rect 315 463 481 481
rect 315 429 333 463
rect 367 429 429 463
rect 463 429 481 463
rect 315 367 481 429
rect 315 333 333 367
rect 367 333 429 367
rect 463 333 481 367
rect 315 315 481 333
<< end >>
