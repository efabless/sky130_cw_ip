magic
tech sky130A
timestamp 1715010268
<< nwell >>
rect 23 35 1253 1063
<< nsubdiff >>
rect 41 1028 94 1045
rect 111 1028 128 1045
rect 145 1028 162 1045
rect 179 1028 196 1045
rect 213 1028 230 1045
rect 247 1028 264 1045
rect 281 1028 298 1045
rect 315 1028 332 1045
rect 349 1028 366 1045
rect 383 1028 400 1045
rect 417 1028 434 1045
rect 451 1028 468 1045
rect 485 1028 502 1045
rect 519 1028 536 1045
rect 553 1028 570 1045
rect 587 1028 604 1045
rect 621 1028 638 1045
rect 655 1028 672 1045
rect 689 1028 706 1045
rect 723 1028 740 1045
rect 757 1028 774 1045
rect 791 1028 808 1045
rect 825 1028 842 1045
rect 859 1028 876 1045
rect 893 1028 910 1045
rect 927 1028 944 1045
rect 961 1028 978 1045
rect 995 1028 1012 1045
rect 1029 1028 1046 1045
rect 1063 1028 1080 1045
rect 1097 1028 1114 1045
rect 1131 1028 1148 1045
rect 1165 1028 1235 1045
rect 41 975 58 1028
rect 41 941 58 958
rect 41 907 58 924
rect 41 873 58 890
rect 41 839 58 856
rect 41 805 58 822
rect 41 771 58 788
rect 41 737 58 754
rect 41 703 58 720
rect 41 669 58 686
rect 41 635 58 652
rect 41 601 58 618
rect 41 567 58 584
rect 41 533 58 550
rect 41 499 58 516
rect 41 465 58 482
rect 41 431 58 448
rect 41 397 58 414
rect 41 363 58 380
rect 41 329 58 346
rect 41 295 58 312
rect 41 261 58 278
rect 41 227 58 244
rect 41 193 58 210
rect 41 159 58 176
rect 41 70 58 142
rect 1218 975 1235 1028
rect 1218 941 1235 958
rect 1218 907 1235 924
rect 1218 873 1235 890
rect 1218 839 1235 856
rect 1218 805 1235 822
rect 1218 771 1235 788
rect 1218 737 1235 754
rect 1218 703 1235 720
rect 1218 669 1235 686
rect 1218 635 1235 652
rect 1218 601 1235 618
rect 1218 567 1235 584
rect 1218 533 1235 550
rect 1218 499 1235 516
rect 1218 465 1235 482
rect 1218 431 1235 448
rect 1218 397 1235 414
rect 1218 363 1235 380
rect 1218 329 1235 346
rect 1218 295 1235 312
rect 1218 261 1235 278
rect 1218 227 1235 244
rect 1218 193 1235 210
rect 1218 159 1235 176
rect 1218 70 1235 142
rect 41 53 128 70
rect 145 53 162 70
rect 179 53 196 70
rect 213 53 230 70
rect 247 53 264 70
rect 281 53 298 70
rect 315 53 332 70
rect 349 53 366 70
rect 383 53 400 70
rect 417 53 434 70
rect 451 53 468 70
rect 485 53 502 70
rect 519 53 536 70
rect 553 53 570 70
rect 587 53 604 70
rect 621 53 638 70
rect 655 53 672 70
rect 689 53 706 70
rect 723 53 740 70
rect 757 53 774 70
rect 791 53 808 70
rect 825 53 842 70
rect 859 53 876 70
rect 893 53 910 70
rect 927 53 944 70
rect 961 53 978 70
rect 995 53 1012 70
rect 1029 53 1046 70
rect 1063 53 1080 70
rect 1097 53 1114 70
rect 1131 53 1148 70
rect 1165 53 1235 70
<< nsubdiffcont >>
rect 94 1028 111 1045
rect 128 1028 145 1045
rect 162 1028 179 1045
rect 196 1028 213 1045
rect 230 1028 247 1045
rect 264 1028 281 1045
rect 298 1028 315 1045
rect 332 1028 349 1045
rect 366 1028 383 1045
rect 400 1028 417 1045
rect 434 1028 451 1045
rect 468 1028 485 1045
rect 502 1028 519 1045
rect 536 1028 553 1045
rect 570 1028 587 1045
rect 604 1028 621 1045
rect 638 1028 655 1045
rect 672 1028 689 1045
rect 706 1028 723 1045
rect 740 1028 757 1045
rect 774 1028 791 1045
rect 808 1028 825 1045
rect 842 1028 859 1045
rect 876 1028 893 1045
rect 910 1028 927 1045
rect 944 1028 961 1045
rect 978 1028 995 1045
rect 1012 1028 1029 1045
rect 1046 1028 1063 1045
rect 1080 1028 1097 1045
rect 1114 1028 1131 1045
rect 1148 1028 1165 1045
rect 41 958 58 975
rect 41 924 58 941
rect 41 890 58 907
rect 41 856 58 873
rect 41 822 58 839
rect 41 788 58 805
rect 41 754 58 771
rect 41 720 58 737
rect 41 686 58 703
rect 41 652 58 669
rect 41 618 58 635
rect 41 584 58 601
rect 41 550 58 567
rect 41 516 58 533
rect 41 482 58 499
rect 41 448 58 465
rect 41 414 58 431
rect 41 380 58 397
rect 41 346 58 363
rect 41 312 58 329
rect 41 278 58 295
rect 41 244 58 261
rect 41 210 58 227
rect 41 176 58 193
rect 41 142 58 159
rect 1218 958 1235 975
rect 1218 924 1235 941
rect 1218 890 1235 907
rect 1218 856 1235 873
rect 1218 822 1235 839
rect 1218 788 1235 805
rect 1218 754 1235 771
rect 1218 720 1235 737
rect 1218 686 1235 703
rect 1218 652 1235 669
rect 1218 618 1235 635
rect 1218 584 1235 601
rect 1218 550 1235 567
rect 1218 516 1235 533
rect 1218 482 1235 499
rect 1218 448 1235 465
rect 1218 414 1235 431
rect 1218 380 1235 397
rect 1218 346 1235 363
rect 1218 312 1235 329
rect 1218 278 1235 295
rect 1218 244 1235 261
rect 1218 210 1235 227
rect 1218 176 1235 193
rect 1218 142 1235 159
rect 128 53 145 70
rect 162 53 179 70
rect 196 53 213 70
rect 230 53 247 70
rect 264 53 281 70
rect 298 53 315 70
rect 332 53 349 70
rect 366 53 383 70
rect 400 53 417 70
rect 434 53 451 70
rect 468 53 485 70
rect 502 53 519 70
rect 536 53 553 70
rect 570 53 587 70
rect 604 53 621 70
rect 638 53 655 70
rect 672 53 689 70
rect 706 53 723 70
rect 740 53 757 70
rect 774 53 791 70
rect 808 53 825 70
rect 842 53 859 70
rect 876 53 893 70
rect 910 53 927 70
rect 944 53 961 70
rect 978 53 995 70
rect 1012 53 1029 70
rect 1046 53 1063 70
rect 1080 53 1097 70
rect 1114 53 1131 70
rect 1148 53 1165 70
<< locali >>
rect 41 1028 94 1045
rect 111 1028 128 1045
rect 145 1028 162 1045
rect 179 1028 196 1045
rect 213 1028 230 1045
rect 247 1028 264 1045
rect 281 1028 298 1045
rect 315 1028 332 1045
rect 349 1028 366 1045
rect 383 1028 400 1045
rect 417 1028 434 1045
rect 451 1028 468 1045
rect 485 1028 502 1045
rect 519 1028 536 1045
rect 553 1028 570 1045
rect 587 1028 604 1045
rect 621 1028 638 1045
rect 655 1028 672 1045
rect 689 1028 706 1045
rect 723 1028 740 1045
rect 757 1028 774 1045
rect 791 1028 808 1045
rect 825 1028 842 1045
rect 859 1028 876 1045
rect 893 1028 910 1045
rect 927 1028 944 1045
rect 961 1028 978 1045
rect 995 1028 1012 1045
rect 1029 1028 1046 1045
rect 1063 1028 1080 1045
rect 1097 1028 1114 1045
rect 1131 1028 1148 1045
rect 1165 1028 1235 1045
rect 41 975 58 1028
rect 41 941 58 958
rect 41 907 58 924
rect 41 873 58 890
rect 41 839 58 856
rect 41 805 58 822
rect 41 771 58 788
rect 41 737 58 754
rect 41 703 58 720
rect 41 669 58 686
rect 41 635 58 652
rect 41 601 58 618
rect 41 567 58 584
rect 41 533 58 550
rect 41 499 58 516
rect 41 465 58 482
rect 41 431 58 448
rect 41 397 58 414
rect 41 363 58 380
rect 41 329 58 346
rect 41 295 58 312
rect 41 261 58 278
rect 41 227 58 244
rect 41 193 58 210
rect 41 159 58 176
rect 41 70 58 142
rect 1218 975 1235 1028
rect 1218 941 1235 958
rect 1218 907 1235 924
rect 1218 873 1235 890
rect 1218 839 1235 856
rect 1218 805 1235 822
rect 1218 771 1235 788
rect 1218 737 1235 754
rect 1218 703 1235 720
rect 1218 669 1235 686
rect 1218 635 1235 652
rect 1218 601 1235 618
rect 1218 567 1235 584
rect 1218 533 1235 550
rect 1218 499 1235 516
rect 1218 465 1235 482
rect 1218 431 1235 448
rect 1218 397 1235 414
rect 1218 363 1235 380
rect 1218 329 1235 346
rect 1218 295 1235 312
rect 1218 261 1235 278
rect 1218 227 1235 244
rect 1218 193 1235 210
rect 1218 159 1235 176
rect 1218 70 1235 142
rect 41 53 128 70
rect 145 53 162 70
rect 179 53 196 70
rect 213 53 230 70
rect 247 53 264 70
rect 281 53 298 70
rect 315 53 332 70
rect 349 53 366 70
rect 383 53 400 70
rect 417 53 434 70
rect 451 53 468 70
rect 485 53 502 70
rect 519 53 536 70
rect 553 53 570 70
rect 587 53 604 70
rect 621 53 638 70
rect 655 53 672 70
rect 689 53 706 70
rect 723 53 740 70
rect 757 53 774 70
rect 791 53 808 70
rect 825 53 842 70
rect 859 53 876 70
rect 893 53 910 70
rect 927 53 944 70
rect 961 53 978 70
rect 995 53 1012 70
rect 1029 53 1046 70
rect 1063 53 1080 70
rect 1097 53 1114 70
rect 1131 53 1148 70
rect 1165 53 1235 70
<< properties >>
string path 1.150 51.825 61.325 51.825 61.325 3.075 2.475 3.075 2.475 51.825 
<< end >>
