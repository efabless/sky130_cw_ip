magic
tech sky130A
magscale 1 2
timestamp 1715010268
<< pwell >>
rect 735 4326 1393 4412
rect 735 3911 821 4326
rect 1307 3911 1393 4326
rect 735 3825 1393 3911
<< psubdiff >>
rect 761 4352 929 4386
rect 963 4352 997 4386
rect 1031 4352 1065 4386
rect 1099 4352 1133 4386
rect 1167 4352 1367 4386
rect 761 4186 795 4352
rect 761 4118 795 4152
rect 761 3885 795 4084
rect 1333 4186 1367 4352
rect 1333 4118 1367 4152
rect 1333 3885 1367 4084
rect 761 3851 997 3885
rect 1031 3851 1065 3885
rect 1099 3851 1133 3885
rect 1167 3851 1367 3885
<< psubdiffcont >>
rect 929 4352 963 4386
rect 997 4352 1031 4386
rect 1065 4352 1099 4386
rect 1133 4352 1167 4386
rect 761 4152 795 4186
rect 761 4084 795 4118
rect 1333 4152 1367 4186
rect 1333 4084 1367 4118
rect 997 3851 1031 3885
rect 1065 3851 1099 3885
rect 1133 3851 1167 3885
<< locali >>
rect 761 4352 929 4386
rect 963 4352 997 4386
rect 1031 4352 1065 4386
rect 1099 4352 1133 4386
rect 1167 4352 1367 4386
rect 761 4186 795 4352
rect 761 4118 795 4152
rect 761 3885 795 4084
rect 1333 4186 1367 4352
rect 1333 4118 1367 4152
rect 1333 3885 1367 4084
rect 761 3851 997 3885
rect 1031 3851 1065 3885
rect 1099 3851 1133 3885
rect 1167 3851 1367 3885
<< properties >>
string path 18.400 109.225 33.750 109.225 33.750 96.700 19.450 96.700 19.450 109.225 
<< end >>
