magic
tech sky130A
magscale 1 2
timestamp 1715615611
<< pwell >>
rect 407 3153 2959 3239
rect 407 395 2872 3153
rect 2873 395 2959 3153
rect 407 309 2959 395
<< psubdiff >>
rect 433 3179 591 3213
rect 625 3179 659 3213
rect 693 3179 727 3213
rect 761 3179 795 3213
rect 829 3179 863 3213
rect 897 3179 931 3213
rect 965 3179 999 3213
rect 1033 3179 1067 3213
rect 1101 3179 1135 3213
rect 1169 3179 1203 3213
rect 1237 3179 1271 3213
rect 1305 3179 1339 3213
rect 1373 3179 1407 3213
rect 1441 3179 1475 3213
rect 1509 3179 1543 3213
rect 1577 3179 1611 3213
rect 1645 3179 1679 3213
rect 1713 3179 1747 3213
rect 1781 3179 1815 3213
rect 1849 3179 1883 3213
rect 1917 3179 1951 3213
rect 1985 3179 2019 3213
rect 2053 3179 2087 3213
rect 2121 3179 2155 3213
rect 2189 3179 2223 3213
rect 2257 3179 2291 3213
rect 2325 3179 2359 3213
rect 2393 3179 2427 3213
rect 2461 3179 2495 3213
rect 2529 3179 2563 3213
rect 2597 3179 2631 3213
rect 2665 3179 2699 3213
rect 2733 3179 2933 3213
rect 433 2962 467 3179
rect 433 2894 467 2928
rect 433 2826 467 2860
rect 433 2758 467 2792
rect 433 2690 467 2724
rect 433 2622 467 2656
rect 433 2554 467 2588
rect 433 2486 467 2520
rect 433 2418 467 2452
rect 433 2350 467 2384
rect 433 2282 467 2316
rect 433 2214 467 2248
rect 433 2146 467 2180
rect 433 2078 467 2112
rect 433 2010 467 2044
rect 433 1942 467 1976
rect 433 1874 467 1908
rect 433 1806 467 1840
rect 433 1738 467 1772
rect 433 1670 467 1704
rect 433 1602 467 1636
rect 433 1534 467 1568
rect 433 1466 467 1500
rect 433 1398 467 1432
rect 433 1330 467 1364
rect 433 1262 467 1296
rect 433 1194 467 1228
rect 433 1126 467 1160
rect 433 1058 467 1092
rect 433 990 467 1024
rect 433 922 467 956
rect 433 854 467 888
rect 433 786 467 820
rect 433 718 467 752
rect 433 650 467 684
rect 433 582 467 616
rect 433 369 467 548
rect 2899 2962 2933 3179
rect 2899 2894 2933 2928
rect 2899 2826 2933 2860
rect 2899 2758 2933 2792
rect 2899 2690 2933 2724
rect 2899 2622 2933 2656
rect 2899 2554 2933 2588
rect 2899 2486 2933 2520
rect 2899 2418 2933 2452
rect 2899 2350 2933 2384
rect 2899 2282 2933 2316
rect 2899 2214 2933 2248
rect 2899 2146 2933 2180
rect 2899 2078 2933 2112
rect 2899 2010 2933 2044
rect 2899 1942 2933 1976
rect 2899 1874 2933 1908
rect 2899 1806 2933 1840
rect 2899 1738 2933 1772
rect 2899 1670 2933 1704
rect 2899 1602 2933 1636
rect 2899 1534 2933 1568
rect 2899 1466 2933 1500
rect 2899 1398 2933 1432
rect 2899 1330 2933 1364
rect 2899 1262 2933 1296
rect 2899 1194 2933 1228
rect 2899 1126 2933 1160
rect 2899 1058 2933 1092
rect 2899 990 2933 1024
rect 2899 922 2933 956
rect 2899 854 2933 888
rect 2899 786 2933 820
rect 2899 718 2933 752
rect 2899 650 2933 684
rect 2899 582 2933 616
rect 2899 369 2933 548
rect 433 335 659 369
rect 693 335 727 369
rect 761 335 795 369
rect 829 335 863 369
rect 897 335 931 369
rect 965 335 999 369
rect 1033 335 1067 369
rect 1101 335 1135 369
rect 1169 335 1203 369
rect 1237 335 1271 369
rect 1305 335 1339 369
rect 1373 335 1407 369
rect 1441 335 1475 369
rect 1509 335 1543 369
rect 1577 335 1611 369
rect 1645 335 1679 369
rect 1713 335 1747 369
rect 1781 335 1815 369
rect 1849 335 1883 369
rect 1917 335 1951 369
rect 1985 335 2019 369
rect 2053 335 2087 369
rect 2121 335 2155 369
rect 2189 335 2223 369
rect 2257 335 2291 369
rect 2325 335 2359 369
rect 2393 335 2427 369
rect 2461 335 2495 369
rect 2529 335 2563 369
rect 2597 335 2631 369
rect 2665 335 2699 369
rect 2733 335 2933 369
<< psubdiffcont >>
rect 591 3179 625 3213
rect 659 3179 693 3213
rect 727 3179 761 3213
rect 795 3179 829 3213
rect 863 3179 897 3213
rect 931 3179 965 3213
rect 999 3179 1033 3213
rect 1067 3179 1101 3213
rect 1135 3179 1169 3213
rect 1203 3179 1237 3213
rect 1271 3179 1305 3213
rect 1339 3179 1373 3213
rect 1407 3179 1441 3213
rect 1475 3179 1509 3213
rect 1543 3179 1577 3213
rect 1611 3179 1645 3213
rect 1679 3179 1713 3213
rect 1747 3179 1781 3213
rect 1815 3179 1849 3213
rect 1883 3179 1917 3213
rect 1951 3179 1985 3213
rect 2019 3179 2053 3213
rect 2087 3179 2121 3213
rect 2155 3179 2189 3213
rect 2223 3179 2257 3213
rect 2291 3179 2325 3213
rect 2359 3179 2393 3213
rect 2427 3179 2461 3213
rect 2495 3179 2529 3213
rect 2563 3179 2597 3213
rect 2631 3179 2665 3213
rect 2699 3179 2733 3213
rect 433 2928 467 2962
rect 433 2860 467 2894
rect 433 2792 467 2826
rect 433 2724 467 2758
rect 433 2656 467 2690
rect 433 2588 467 2622
rect 433 2520 467 2554
rect 433 2452 467 2486
rect 433 2384 467 2418
rect 433 2316 467 2350
rect 433 2248 467 2282
rect 433 2180 467 2214
rect 433 2112 467 2146
rect 433 2044 467 2078
rect 433 1976 467 2010
rect 433 1908 467 1942
rect 433 1840 467 1874
rect 433 1772 467 1806
rect 433 1704 467 1738
rect 433 1636 467 1670
rect 433 1568 467 1602
rect 433 1500 467 1534
rect 433 1432 467 1466
rect 433 1364 467 1398
rect 433 1296 467 1330
rect 433 1228 467 1262
rect 433 1160 467 1194
rect 433 1092 467 1126
rect 433 1024 467 1058
rect 433 956 467 990
rect 433 888 467 922
rect 433 820 467 854
rect 433 752 467 786
rect 433 684 467 718
rect 433 616 467 650
rect 433 548 467 582
rect 2899 2928 2933 2962
rect 2899 2860 2933 2894
rect 2899 2792 2933 2826
rect 2899 2724 2933 2758
rect 2899 2656 2933 2690
rect 2899 2588 2933 2622
rect 2899 2520 2933 2554
rect 2899 2452 2933 2486
rect 2899 2384 2933 2418
rect 2899 2316 2933 2350
rect 2899 2248 2933 2282
rect 2899 2180 2933 2214
rect 2899 2112 2933 2146
rect 2899 2044 2933 2078
rect 2899 1976 2933 2010
rect 2899 1908 2933 1942
rect 2899 1840 2933 1874
rect 2899 1772 2933 1806
rect 2899 1704 2933 1738
rect 2899 1636 2933 1670
rect 2899 1568 2933 1602
rect 2899 1500 2933 1534
rect 2899 1432 2933 1466
rect 2899 1364 2933 1398
rect 2899 1296 2933 1330
rect 2899 1228 2933 1262
rect 2899 1160 2933 1194
rect 2899 1092 2933 1126
rect 2899 1024 2933 1058
rect 2899 956 2933 990
rect 2899 888 2933 922
rect 2899 820 2933 854
rect 2899 752 2933 786
rect 2899 684 2933 718
rect 2899 616 2933 650
rect 2899 548 2933 582
rect 659 335 693 369
rect 727 335 761 369
rect 795 335 829 369
rect 863 335 897 369
rect 931 335 965 369
rect 999 335 1033 369
rect 1067 335 1101 369
rect 1135 335 1169 369
rect 1203 335 1237 369
rect 1271 335 1305 369
rect 1339 335 1373 369
rect 1407 335 1441 369
rect 1475 335 1509 369
rect 1543 335 1577 369
rect 1611 335 1645 369
rect 1679 335 1713 369
rect 1747 335 1781 369
rect 1815 335 1849 369
rect 1883 335 1917 369
rect 1951 335 1985 369
rect 2019 335 2053 369
rect 2087 335 2121 369
rect 2155 335 2189 369
rect 2223 335 2257 369
rect 2291 335 2325 369
rect 2359 335 2393 369
rect 2427 335 2461 369
rect 2495 335 2529 369
rect 2563 335 2597 369
rect 2631 335 2665 369
rect 2699 335 2733 369
<< locali >>
rect 433 3179 591 3213
rect 625 3179 659 3213
rect 693 3179 727 3213
rect 761 3179 795 3213
rect 829 3179 863 3213
rect 897 3179 931 3213
rect 965 3179 999 3213
rect 1033 3179 1067 3213
rect 1101 3179 1135 3213
rect 1169 3179 1203 3213
rect 1237 3179 1271 3213
rect 1305 3179 1339 3213
rect 1373 3179 1407 3213
rect 1441 3179 1475 3213
rect 1509 3179 1543 3213
rect 1577 3179 1611 3213
rect 1645 3179 1679 3213
rect 1713 3179 1747 3213
rect 1781 3179 1815 3213
rect 1849 3179 1883 3213
rect 1917 3179 1951 3213
rect 1985 3179 2019 3213
rect 2053 3179 2087 3213
rect 2121 3179 2155 3213
rect 2189 3179 2223 3213
rect 2257 3179 2291 3213
rect 2325 3179 2359 3213
rect 2393 3179 2427 3213
rect 2461 3179 2495 3213
rect 2529 3179 2563 3213
rect 2597 3179 2631 3213
rect 2665 3179 2699 3213
rect 2733 3179 2933 3213
rect 433 2962 467 3179
rect 433 2894 467 2928
rect 433 2826 467 2860
rect 433 2758 467 2792
rect 433 2690 467 2724
rect 433 2622 467 2656
rect 433 2554 467 2588
rect 433 2486 467 2520
rect 433 2418 467 2452
rect 433 2350 467 2384
rect 433 2282 467 2316
rect 433 2214 467 2248
rect 433 2146 467 2180
rect 433 2078 467 2112
rect 433 2010 467 2044
rect 433 1942 467 1976
rect 433 1874 467 1908
rect 433 1806 467 1840
rect 433 1738 467 1772
rect 433 1670 467 1704
rect 433 1602 467 1636
rect 433 1534 467 1568
rect 433 1466 467 1500
rect 433 1398 467 1432
rect 433 1330 467 1364
rect 433 1262 467 1296
rect 433 1194 467 1228
rect 433 1126 467 1160
rect 433 1058 467 1092
rect 433 990 467 1024
rect 433 922 467 956
rect 433 854 467 888
rect 433 786 467 820
rect 433 718 467 752
rect 433 650 467 684
rect 433 582 467 616
rect 433 369 467 548
rect 2899 2962 2933 3179
rect 2899 2894 2933 2928
rect 2899 2826 2933 2860
rect 2899 2758 2933 2792
rect 2899 2690 2933 2724
rect 2899 2622 2933 2656
rect 2899 2554 2933 2588
rect 2899 2486 2933 2520
rect 2899 2418 2933 2452
rect 2899 2350 2933 2384
rect 2899 2282 2933 2316
rect 2899 2214 2933 2248
rect 2899 2146 2933 2180
rect 2899 2078 2933 2112
rect 2899 2010 2933 2044
rect 2899 1942 2933 1976
rect 2899 1874 2933 1908
rect 2899 1806 2933 1840
rect 2899 1738 2933 1772
rect 2899 1670 2933 1704
rect 2899 1602 2933 1636
rect 2899 1534 2933 1568
rect 2899 1466 2933 1500
rect 2899 1398 2933 1432
rect 2899 1330 2933 1364
rect 2899 1262 2933 1296
rect 2899 1194 2933 1228
rect 2899 1126 2933 1160
rect 2899 1058 2933 1092
rect 2899 990 2933 1024
rect 2899 922 2933 956
rect 2899 854 2933 888
rect 2899 786 2933 820
rect 2899 718 2933 752
rect 2899 650 2933 684
rect 2899 582 2933 616
rect 2899 369 2933 548
rect 433 335 659 369
rect 693 335 727 369
rect 761 335 795 369
rect 829 335 863 369
rect 897 335 931 369
rect 965 335 999 369
rect 1033 335 1067 369
rect 1101 335 1135 369
rect 1169 335 1203 369
rect 1237 335 1271 369
rect 1305 335 1339 369
rect 1373 335 1407 369
rect 1441 335 1475 369
rect 1509 335 1543 369
rect 1577 335 1611 369
rect 1645 335 1679 369
rect 1713 335 1747 369
rect 1781 335 1815 369
rect 1849 335 1883 369
rect 1917 335 1951 369
rect 1985 335 2019 369
rect 2053 335 2087 369
rect 2121 335 2155 369
rect 2189 335 2223 369
rect 2257 335 2291 369
rect 2325 335 2359 369
rect 2393 335 2427 369
rect 2461 335 2495 369
rect 2529 335 2563 369
rect 2597 335 2631 369
rect 2665 335 2699 369
rect 2733 335 2933 369
<< properties >>
string path 10.200 79.900 72.900 79.900 72.900 8.800 11.250 8.800 11.250 79.900 
<< end >>
