magic
tech sky130A
magscale 1 2
timestamp 1715625863
<< nwell >>
rect -18157 4978 -7349 8917
<< nsubdiff >>
rect -18121 8847 -18034 8881
rect -18000 8847 -17966 8881
rect -17932 8847 -17898 8881
rect -17864 8847 -17830 8881
rect -17796 8847 -17762 8881
rect -17728 8847 -17694 8881
rect -17660 8847 -17626 8881
rect -17592 8847 -17558 8881
rect -17524 8847 -17490 8881
rect -17456 8847 -17422 8881
rect -17388 8847 -17354 8881
rect -17320 8847 -17286 8881
rect -17252 8847 -17218 8881
rect -17184 8847 -17150 8881
rect -17116 8847 -17082 8881
rect -17048 8847 -17014 8881
rect -16980 8847 -16946 8881
rect -16912 8847 -16878 8881
rect -16844 8847 -16810 8881
rect -16776 8847 -16742 8881
rect -16708 8847 -16674 8881
rect -16640 8847 -16606 8881
rect -16572 8847 -16538 8881
rect -16504 8847 -16470 8881
rect -16436 8847 -16402 8881
rect -16368 8847 -16334 8881
rect -16300 8847 -16266 8881
rect -16232 8847 -16198 8881
rect -16164 8847 -16130 8881
rect -16096 8847 -16062 8881
rect -16028 8847 -15994 8881
rect -15960 8847 -15926 8881
rect -15892 8847 -15858 8881
rect -15824 8847 -15790 8881
rect -15756 8847 -15722 8881
rect -15688 8847 -15654 8881
rect -15620 8847 -15586 8881
rect -15552 8847 -15518 8881
rect -15484 8847 -15450 8881
rect -15416 8847 -15382 8881
rect -15348 8847 -15314 8881
rect -15280 8847 -15246 8881
rect -15212 8847 -15178 8881
rect -15144 8847 -15110 8881
rect -15076 8847 -15042 8881
rect -15008 8847 -14974 8881
rect -14940 8847 -14906 8881
rect -14872 8847 -14838 8881
rect -14804 8847 -14770 8881
rect -14736 8847 -14702 8881
rect -14668 8847 -14634 8881
rect -14600 8847 -14566 8881
rect -14532 8847 -14498 8881
rect -14464 8847 -14430 8881
rect -14396 8847 -14362 8881
rect -14328 8847 -14294 8881
rect -14260 8847 -14226 8881
rect -14192 8847 -14158 8881
rect -14124 8847 -14090 8881
rect -14056 8847 -14022 8881
rect -13988 8847 -13954 8881
rect -13920 8847 -13886 8881
rect -13852 8847 -13818 8881
rect -13784 8847 -13750 8881
rect -13716 8847 -13682 8881
rect -13648 8847 -13614 8881
rect -13580 8847 -13546 8881
rect -13512 8847 -13478 8881
rect -13444 8847 -13410 8881
rect -13376 8847 -13342 8881
rect -13308 8847 -13274 8881
rect -13240 8847 -13206 8881
rect -13172 8847 -13138 8881
rect -13104 8847 -13070 8881
rect -13036 8847 -13002 8881
rect -12968 8847 -12934 8881
rect -12900 8847 -12866 8881
rect -12832 8847 -12798 8881
rect -12764 8847 -12730 8881
rect -12696 8847 -12662 8881
rect -12628 8847 -12594 8881
rect -12560 8847 -12526 8881
rect -12492 8847 -12458 8881
rect -12424 8847 -12390 8881
rect -12356 8847 -12322 8881
rect -12288 8847 -12254 8881
rect -12220 8847 -12186 8881
rect -12152 8847 -12118 8881
rect -12084 8847 -12050 8881
rect -12016 8847 -11982 8881
rect -11948 8847 -11914 8881
rect -11880 8847 -11846 8881
rect -11812 8847 -11778 8881
rect -11744 8847 -11710 8881
rect -11676 8847 -11642 8881
rect -11608 8847 -11574 8881
rect -11540 8847 -11506 8881
rect -11472 8847 -11438 8881
rect -11404 8847 -11370 8881
rect -11336 8847 -11302 8881
rect -11268 8847 -11234 8881
rect -11200 8847 -11166 8881
rect -11132 8847 -11098 8881
rect -11064 8847 -11030 8881
rect -10996 8847 -10962 8881
rect -10928 8847 -10894 8881
rect -10860 8847 -10826 8881
rect -10792 8847 -10758 8881
rect -10724 8847 -10690 8881
rect -10656 8847 -10622 8881
rect -10588 8847 -10554 8881
rect -10520 8847 -10486 8881
rect -10452 8847 -10418 8881
rect -10384 8847 -10350 8881
rect -10316 8847 -10282 8881
rect -10248 8847 -10214 8881
rect -10180 8847 -10146 8881
rect -10112 8847 -10078 8881
rect -10044 8847 -10010 8881
rect -9976 8847 -9942 8881
rect -9908 8847 -9874 8881
rect -9840 8847 -9806 8881
rect -9772 8847 -9738 8881
rect -9704 8847 -9670 8881
rect -9636 8847 -9602 8881
rect -9568 8847 -9534 8881
rect -9500 8847 -9466 8881
rect -9432 8847 -9398 8881
rect -9364 8847 -9330 8881
rect -9296 8847 -9262 8881
rect -9228 8847 -9194 8881
rect -9160 8847 -9126 8881
rect -9092 8847 -9058 8881
rect -9024 8847 -8990 8881
rect -8956 8847 -8922 8881
rect -8888 8847 -8854 8881
rect -8820 8847 -8786 8881
rect -8752 8847 -8718 8881
rect -8684 8847 -8650 8881
rect -8616 8847 -8582 8881
rect -8548 8847 -8514 8881
rect -8480 8847 -8446 8881
rect -8412 8847 -8378 8881
rect -8344 8847 -8310 8881
rect -8276 8847 -8242 8881
rect -8208 8847 -8174 8881
rect -8140 8847 -8106 8881
rect -8072 8847 -8038 8881
rect -8004 8847 -7970 8881
rect -7936 8847 -7902 8881
rect -7868 8847 -7834 8881
rect -7800 8847 -7766 8881
rect -7732 8847 -7698 8881
rect -7664 8847 -7630 8881
rect -7596 8847 -7562 8881
rect -7528 8847 -7385 8881
rect -18121 8741 -18087 8847
rect -18121 8673 -18087 8707
rect -18121 8605 -18087 8639
rect -18121 8537 -18087 8571
rect -18121 8469 -18087 8503
rect -18121 8401 -18087 8435
rect -18121 8333 -18087 8367
rect -18121 8265 -18087 8299
rect -18121 8197 -18087 8231
rect -18121 8129 -18087 8163
rect -18121 8061 -18087 8095
rect -18121 7993 -18087 8027
rect -18121 7925 -18087 7959
rect -18121 7857 -18087 7891
rect -18121 7789 -18087 7823
rect -18121 7721 -18087 7755
rect -18121 7653 -18087 7687
rect -18121 7585 -18087 7619
rect -18121 7517 -18087 7551
rect -18121 7449 -18087 7483
rect -18121 7381 -18087 7415
rect -18121 7313 -18087 7347
rect -18121 7245 -18087 7279
rect -18121 7177 -18087 7211
rect -18121 7109 -18087 7143
rect -18121 7041 -18087 7075
rect -18121 6973 -18087 7007
rect -18121 6905 -18087 6939
rect -18121 6837 -18087 6871
rect -18121 6769 -18087 6803
rect -18121 6701 -18087 6735
rect -18121 6633 -18087 6667
rect -18121 6565 -18087 6599
rect -18121 6497 -18087 6531
rect -18121 6429 -18087 6463
rect -18121 6361 -18087 6395
rect -18121 6293 -18087 6327
rect -18121 6225 -18087 6259
rect -18121 6157 -18087 6191
rect -18121 6089 -18087 6123
rect -18121 6021 -18087 6055
rect -18121 5953 -18087 5987
rect -18121 5885 -18087 5919
rect -18121 5817 -18087 5851
rect -18121 5749 -18087 5783
rect -18121 5681 -18087 5715
rect -18121 5613 -18087 5647
rect -18121 5545 -18087 5579
rect -18121 5477 -18087 5511
rect -18121 5409 -18087 5443
rect -18121 5341 -18087 5375
rect -18121 5273 -18087 5307
rect -18121 5205 -18087 5239
rect -18121 5048 -18087 5171
rect -7419 8741 -7385 8847
rect -7419 8673 -7385 8707
rect -7419 8605 -7385 8639
rect -7419 8537 -7385 8571
rect -7419 8469 -7385 8503
rect -7419 8401 -7385 8435
rect -7419 8333 -7385 8367
rect -7419 8265 -7385 8299
rect -7419 8197 -7385 8231
rect -7419 8129 -7385 8163
rect -7419 8061 -7385 8095
rect -7419 7993 -7385 8027
rect -7419 7925 -7385 7959
rect -7419 7857 -7385 7891
rect -7419 7789 -7385 7823
rect -7419 7721 -7385 7755
rect -7419 7653 -7385 7687
rect -7419 7585 -7385 7619
rect -7419 7517 -7385 7551
rect -7419 7449 -7385 7483
rect -7419 7381 -7385 7415
rect -7419 7313 -7385 7347
rect -7419 7245 -7385 7279
rect -7419 7177 -7385 7211
rect -7419 7109 -7385 7143
rect -7419 7041 -7385 7075
rect -7419 6973 -7385 7007
rect -7419 6905 -7385 6939
rect -7419 6837 -7385 6871
rect -7419 6769 -7385 6803
rect -7419 6701 -7385 6735
rect -7419 6633 -7385 6667
rect -7419 6565 -7385 6599
rect -7419 6497 -7385 6531
rect -7419 6429 -7385 6463
rect -7419 6361 -7385 6395
rect -7419 6293 -7385 6327
rect -7419 6225 -7385 6259
rect -7419 6157 -7385 6191
rect -7419 6089 -7385 6123
rect -7419 6021 -7385 6055
rect -7419 5953 -7385 5987
rect -7419 5885 -7385 5919
rect -7419 5817 -7385 5851
rect -7419 5749 -7385 5783
rect -7419 5681 -7385 5715
rect -7419 5613 -7385 5647
rect -7419 5545 -7385 5579
rect -7419 5477 -7385 5511
rect -7419 5409 -7385 5443
rect -7419 5341 -7385 5375
rect -7419 5273 -7385 5307
rect -7419 5205 -7385 5239
rect -7419 5048 -7385 5171
rect -18121 5014 -17981 5048
rect -17947 5014 -17913 5048
rect -17879 5014 -17845 5048
rect -17811 5014 -17777 5048
rect -17743 5014 -17709 5048
rect -17675 5014 -17641 5048
rect -17607 5014 -17573 5048
rect -17539 5014 -17505 5048
rect -17471 5014 -17437 5048
rect -17403 5014 -17369 5048
rect -17335 5014 -17301 5048
rect -17267 5014 -17233 5048
rect -17199 5014 -17165 5048
rect -17131 5014 -17097 5048
rect -17063 5014 -17029 5048
rect -16995 5014 -16961 5048
rect -16927 5014 -16893 5048
rect -16859 5014 -16825 5048
rect -16791 5014 -16757 5048
rect -16723 5014 -16689 5048
rect -16655 5014 -16621 5048
rect -16587 5014 -16553 5048
rect -16519 5014 -16485 5048
rect -16451 5014 -16417 5048
rect -16383 5014 -16349 5048
rect -16315 5014 -16281 5048
rect -16247 5014 -16213 5048
rect -16179 5014 -16145 5048
rect -16111 5014 -16077 5048
rect -16043 5014 -16009 5048
rect -15975 5014 -15941 5048
rect -15907 5014 -15873 5048
rect -15839 5014 -15805 5048
rect -15771 5014 -15737 5048
rect -15703 5014 -15669 5048
rect -15635 5014 -15601 5048
rect -15567 5014 -15533 5048
rect -15499 5014 -15465 5048
rect -15431 5014 -15397 5048
rect -15363 5014 -15329 5048
rect -15295 5014 -15261 5048
rect -15227 5014 -15193 5048
rect -15159 5014 -15125 5048
rect -15091 5014 -15057 5048
rect -15023 5014 -14989 5048
rect -14955 5014 -14921 5048
rect -14887 5014 -14853 5048
rect -14819 5014 -14785 5048
rect -14751 5014 -14717 5048
rect -14683 5014 -14649 5048
rect -14615 5014 -14581 5048
rect -14547 5014 -14513 5048
rect -14479 5014 -14445 5048
rect -14411 5014 -14377 5048
rect -14343 5014 -14309 5048
rect -14275 5014 -14241 5048
rect -14207 5014 -14173 5048
rect -14139 5014 -14105 5048
rect -14071 5014 -14037 5048
rect -14003 5014 -13969 5048
rect -13935 5014 -13901 5048
rect -13867 5014 -13833 5048
rect -13799 5014 -13765 5048
rect -13731 5014 -13697 5048
rect -13663 5014 -13629 5048
rect -13595 5014 -13561 5048
rect -13527 5014 -13493 5048
rect -13459 5014 -13425 5048
rect -13391 5014 -13357 5048
rect -13323 5014 -13289 5048
rect -13255 5014 -13221 5048
rect -13187 5014 -13153 5048
rect -13119 5014 -13085 5048
rect -13051 5014 -13017 5048
rect -12983 5014 -12949 5048
rect -12915 5014 -12881 5048
rect -12847 5014 -12813 5048
rect -12779 5014 -12745 5048
rect -12711 5014 -12677 5048
rect -12643 5014 -12609 5048
rect -12575 5014 -12541 5048
rect -12507 5014 -12473 5048
rect -12439 5014 -12405 5048
rect -12371 5014 -12337 5048
rect -12303 5014 -12269 5048
rect -12235 5014 -12201 5048
rect -12167 5014 -12133 5048
rect -12099 5014 -12065 5048
rect -12031 5014 -11997 5048
rect -11963 5014 -11929 5048
rect -11895 5014 -11861 5048
rect -11827 5014 -11793 5048
rect -11759 5014 -11725 5048
rect -11691 5014 -11657 5048
rect -11623 5014 -11589 5048
rect -11555 5014 -11521 5048
rect -11487 5014 -11453 5048
rect -11419 5014 -11385 5048
rect -11351 5014 -11317 5048
rect -11283 5014 -11249 5048
rect -11215 5014 -11181 5048
rect -11147 5014 -11113 5048
rect -11079 5014 -11045 5048
rect -11011 5014 -10977 5048
rect -10943 5014 -10909 5048
rect -10875 5014 -10841 5048
rect -10807 5014 -10773 5048
rect -10739 5014 -10705 5048
rect -10671 5014 -10637 5048
rect -10603 5014 -10569 5048
rect -10535 5014 -10501 5048
rect -10467 5014 -10433 5048
rect -10399 5014 -10365 5048
rect -10331 5014 -10297 5048
rect -10263 5014 -10229 5048
rect -10195 5014 -10161 5048
rect -10127 5014 -10093 5048
rect -10059 5014 -10025 5048
rect -9991 5014 -9957 5048
rect -9923 5014 -9889 5048
rect -9855 5014 -9821 5048
rect -9787 5014 -9753 5048
rect -9719 5014 -9685 5048
rect -9651 5014 -9617 5048
rect -9583 5014 -9549 5048
rect -9515 5014 -9481 5048
rect -9447 5014 -9413 5048
rect -9379 5014 -9345 5048
rect -9311 5014 -9277 5048
rect -9243 5014 -9209 5048
rect -9175 5014 -9141 5048
rect -9107 5014 -9073 5048
rect -9039 5014 -9005 5048
rect -8971 5014 -8937 5048
rect -8903 5014 -8869 5048
rect -8835 5014 -8801 5048
rect -8767 5014 -8733 5048
rect -8699 5014 -8665 5048
rect -8631 5014 -8597 5048
rect -8563 5014 -8529 5048
rect -8495 5014 -8461 5048
rect -8427 5014 -8393 5048
rect -8359 5014 -8325 5048
rect -8291 5014 -8257 5048
rect -8223 5014 -8189 5048
rect -8155 5014 -8121 5048
rect -8087 5014 -8053 5048
rect -8019 5014 -7985 5048
rect -7951 5014 -7917 5048
rect -7883 5014 -7849 5048
rect -7815 5014 -7781 5048
rect -7747 5014 -7713 5048
rect -7679 5014 -7645 5048
rect -7611 5014 -7577 5048
rect -7543 5014 -7385 5048
<< nsubdiffcont >>
rect -18034 8847 -18000 8881
rect -17966 8847 -17932 8881
rect -17898 8847 -17864 8881
rect -17830 8847 -17796 8881
rect -17762 8847 -17728 8881
rect -17694 8847 -17660 8881
rect -17626 8847 -17592 8881
rect -17558 8847 -17524 8881
rect -17490 8847 -17456 8881
rect -17422 8847 -17388 8881
rect -17354 8847 -17320 8881
rect -17286 8847 -17252 8881
rect -17218 8847 -17184 8881
rect -17150 8847 -17116 8881
rect -17082 8847 -17048 8881
rect -17014 8847 -16980 8881
rect -16946 8847 -16912 8881
rect -16878 8847 -16844 8881
rect -16810 8847 -16776 8881
rect -16742 8847 -16708 8881
rect -16674 8847 -16640 8881
rect -16606 8847 -16572 8881
rect -16538 8847 -16504 8881
rect -16470 8847 -16436 8881
rect -16402 8847 -16368 8881
rect -16334 8847 -16300 8881
rect -16266 8847 -16232 8881
rect -16198 8847 -16164 8881
rect -16130 8847 -16096 8881
rect -16062 8847 -16028 8881
rect -15994 8847 -15960 8881
rect -15926 8847 -15892 8881
rect -15858 8847 -15824 8881
rect -15790 8847 -15756 8881
rect -15722 8847 -15688 8881
rect -15654 8847 -15620 8881
rect -15586 8847 -15552 8881
rect -15518 8847 -15484 8881
rect -15450 8847 -15416 8881
rect -15382 8847 -15348 8881
rect -15314 8847 -15280 8881
rect -15246 8847 -15212 8881
rect -15178 8847 -15144 8881
rect -15110 8847 -15076 8881
rect -15042 8847 -15008 8881
rect -14974 8847 -14940 8881
rect -14906 8847 -14872 8881
rect -14838 8847 -14804 8881
rect -14770 8847 -14736 8881
rect -14702 8847 -14668 8881
rect -14634 8847 -14600 8881
rect -14566 8847 -14532 8881
rect -14498 8847 -14464 8881
rect -14430 8847 -14396 8881
rect -14362 8847 -14328 8881
rect -14294 8847 -14260 8881
rect -14226 8847 -14192 8881
rect -14158 8847 -14124 8881
rect -14090 8847 -14056 8881
rect -14022 8847 -13988 8881
rect -13954 8847 -13920 8881
rect -13886 8847 -13852 8881
rect -13818 8847 -13784 8881
rect -13750 8847 -13716 8881
rect -13682 8847 -13648 8881
rect -13614 8847 -13580 8881
rect -13546 8847 -13512 8881
rect -13478 8847 -13444 8881
rect -13410 8847 -13376 8881
rect -13342 8847 -13308 8881
rect -13274 8847 -13240 8881
rect -13206 8847 -13172 8881
rect -13138 8847 -13104 8881
rect -13070 8847 -13036 8881
rect -13002 8847 -12968 8881
rect -12934 8847 -12900 8881
rect -12866 8847 -12832 8881
rect -12798 8847 -12764 8881
rect -12730 8847 -12696 8881
rect -12662 8847 -12628 8881
rect -12594 8847 -12560 8881
rect -12526 8847 -12492 8881
rect -12458 8847 -12424 8881
rect -12390 8847 -12356 8881
rect -12322 8847 -12288 8881
rect -12254 8847 -12220 8881
rect -12186 8847 -12152 8881
rect -12118 8847 -12084 8881
rect -12050 8847 -12016 8881
rect -11982 8847 -11948 8881
rect -11914 8847 -11880 8881
rect -11846 8847 -11812 8881
rect -11778 8847 -11744 8881
rect -11710 8847 -11676 8881
rect -11642 8847 -11608 8881
rect -11574 8847 -11540 8881
rect -11506 8847 -11472 8881
rect -11438 8847 -11404 8881
rect -11370 8847 -11336 8881
rect -11302 8847 -11268 8881
rect -11234 8847 -11200 8881
rect -11166 8847 -11132 8881
rect -11098 8847 -11064 8881
rect -11030 8847 -10996 8881
rect -10962 8847 -10928 8881
rect -10894 8847 -10860 8881
rect -10826 8847 -10792 8881
rect -10758 8847 -10724 8881
rect -10690 8847 -10656 8881
rect -10622 8847 -10588 8881
rect -10554 8847 -10520 8881
rect -10486 8847 -10452 8881
rect -10418 8847 -10384 8881
rect -10350 8847 -10316 8881
rect -10282 8847 -10248 8881
rect -10214 8847 -10180 8881
rect -10146 8847 -10112 8881
rect -10078 8847 -10044 8881
rect -10010 8847 -9976 8881
rect -9942 8847 -9908 8881
rect -9874 8847 -9840 8881
rect -9806 8847 -9772 8881
rect -9738 8847 -9704 8881
rect -9670 8847 -9636 8881
rect -9602 8847 -9568 8881
rect -9534 8847 -9500 8881
rect -9466 8847 -9432 8881
rect -9398 8847 -9364 8881
rect -9330 8847 -9296 8881
rect -9262 8847 -9228 8881
rect -9194 8847 -9160 8881
rect -9126 8847 -9092 8881
rect -9058 8847 -9024 8881
rect -8990 8847 -8956 8881
rect -8922 8847 -8888 8881
rect -8854 8847 -8820 8881
rect -8786 8847 -8752 8881
rect -8718 8847 -8684 8881
rect -8650 8847 -8616 8881
rect -8582 8847 -8548 8881
rect -8514 8847 -8480 8881
rect -8446 8847 -8412 8881
rect -8378 8847 -8344 8881
rect -8310 8847 -8276 8881
rect -8242 8847 -8208 8881
rect -8174 8847 -8140 8881
rect -8106 8847 -8072 8881
rect -8038 8847 -8004 8881
rect -7970 8847 -7936 8881
rect -7902 8847 -7868 8881
rect -7834 8847 -7800 8881
rect -7766 8847 -7732 8881
rect -7698 8847 -7664 8881
rect -7630 8847 -7596 8881
rect -7562 8847 -7528 8881
rect -18121 8707 -18087 8741
rect -18121 8639 -18087 8673
rect -18121 8571 -18087 8605
rect -18121 8503 -18087 8537
rect -18121 8435 -18087 8469
rect -18121 8367 -18087 8401
rect -18121 8299 -18087 8333
rect -18121 8231 -18087 8265
rect -18121 8163 -18087 8197
rect -18121 8095 -18087 8129
rect -18121 8027 -18087 8061
rect -18121 7959 -18087 7993
rect -18121 7891 -18087 7925
rect -18121 7823 -18087 7857
rect -18121 7755 -18087 7789
rect -18121 7687 -18087 7721
rect -18121 7619 -18087 7653
rect -18121 7551 -18087 7585
rect -18121 7483 -18087 7517
rect -18121 7415 -18087 7449
rect -18121 7347 -18087 7381
rect -18121 7279 -18087 7313
rect -18121 7211 -18087 7245
rect -18121 7143 -18087 7177
rect -18121 7075 -18087 7109
rect -18121 7007 -18087 7041
rect -18121 6939 -18087 6973
rect -18121 6871 -18087 6905
rect -18121 6803 -18087 6837
rect -18121 6735 -18087 6769
rect -18121 6667 -18087 6701
rect -18121 6599 -18087 6633
rect -18121 6531 -18087 6565
rect -18121 6463 -18087 6497
rect -18121 6395 -18087 6429
rect -18121 6327 -18087 6361
rect -18121 6259 -18087 6293
rect -18121 6191 -18087 6225
rect -18121 6123 -18087 6157
rect -18121 6055 -18087 6089
rect -18121 5987 -18087 6021
rect -18121 5919 -18087 5953
rect -18121 5851 -18087 5885
rect -18121 5783 -18087 5817
rect -18121 5715 -18087 5749
rect -18121 5647 -18087 5681
rect -18121 5579 -18087 5613
rect -18121 5511 -18087 5545
rect -18121 5443 -18087 5477
rect -18121 5375 -18087 5409
rect -18121 5307 -18087 5341
rect -18121 5239 -18087 5273
rect -18121 5171 -18087 5205
rect -7419 8707 -7385 8741
rect -7419 8639 -7385 8673
rect -7419 8571 -7385 8605
rect -7419 8503 -7385 8537
rect -7419 8435 -7385 8469
rect -7419 8367 -7385 8401
rect -7419 8299 -7385 8333
rect -7419 8231 -7385 8265
rect -7419 8163 -7385 8197
rect -7419 8095 -7385 8129
rect -7419 8027 -7385 8061
rect -7419 7959 -7385 7993
rect -7419 7891 -7385 7925
rect -7419 7823 -7385 7857
rect -7419 7755 -7385 7789
rect -7419 7687 -7385 7721
rect -7419 7619 -7385 7653
rect -7419 7551 -7385 7585
rect -7419 7483 -7385 7517
rect -7419 7415 -7385 7449
rect -7419 7347 -7385 7381
rect -7419 7279 -7385 7313
rect -7419 7211 -7385 7245
rect -7419 7143 -7385 7177
rect -7419 7075 -7385 7109
rect -7419 7007 -7385 7041
rect -7419 6939 -7385 6973
rect -7419 6871 -7385 6905
rect -7419 6803 -7385 6837
rect -7419 6735 -7385 6769
rect -7419 6667 -7385 6701
rect -7419 6599 -7385 6633
rect -7419 6531 -7385 6565
rect -7419 6463 -7385 6497
rect -7419 6395 -7385 6429
rect -7419 6327 -7385 6361
rect -7419 6259 -7385 6293
rect -7419 6191 -7385 6225
rect -7419 6123 -7385 6157
rect -7419 6055 -7385 6089
rect -7419 5987 -7385 6021
rect -7419 5919 -7385 5953
rect -7419 5851 -7385 5885
rect -7419 5783 -7385 5817
rect -7419 5715 -7385 5749
rect -7419 5647 -7385 5681
rect -7419 5579 -7385 5613
rect -7419 5511 -7385 5545
rect -7419 5443 -7385 5477
rect -7419 5375 -7385 5409
rect -7419 5307 -7385 5341
rect -7419 5239 -7385 5273
rect -7419 5171 -7385 5205
rect -17981 5014 -17947 5048
rect -17913 5014 -17879 5048
rect -17845 5014 -17811 5048
rect -17777 5014 -17743 5048
rect -17709 5014 -17675 5048
rect -17641 5014 -17607 5048
rect -17573 5014 -17539 5048
rect -17505 5014 -17471 5048
rect -17437 5014 -17403 5048
rect -17369 5014 -17335 5048
rect -17301 5014 -17267 5048
rect -17233 5014 -17199 5048
rect -17165 5014 -17131 5048
rect -17097 5014 -17063 5048
rect -17029 5014 -16995 5048
rect -16961 5014 -16927 5048
rect -16893 5014 -16859 5048
rect -16825 5014 -16791 5048
rect -16757 5014 -16723 5048
rect -16689 5014 -16655 5048
rect -16621 5014 -16587 5048
rect -16553 5014 -16519 5048
rect -16485 5014 -16451 5048
rect -16417 5014 -16383 5048
rect -16349 5014 -16315 5048
rect -16281 5014 -16247 5048
rect -16213 5014 -16179 5048
rect -16145 5014 -16111 5048
rect -16077 5014 -16043 5048
rect -16009 5014 -15975 5048
rect -15941 5014 -15907 5048
rect -15873 5014 -15839 5048
rect -15805 5014 -15771 5048
rect -15737 5014 -15703 5048
rect -15669 5014 -15635 5048
rect -15601 5014 -15567 5048
rect -15533 5014 -15499 5048
rect -15465 5014 -15431 5048
rect -15397 5014 -15363 5048
rect -15329 5014 -15295 5048
rect -15261 5014 -15227 5048
rect -15193 5014 -15159 5048
rect -15125 5014 -15091 5048
rect -15057 5014 -15023 5048
rect -14989 5014 -14955 5048
rect -14921 5014 -14887 5048
rect -14853 5014 -14819 5048
rect -14785 5014 -14751 5048
rect -14717 5014 -14683 5048
rect -14649 5014 -14615 5048
rect -14581 5014 -14547 5048
rect -14513 5014 -14479 5048
rect -14445 5014 -14411 5048
rect -14377 5014 -14343 5048
rect -14309 5014 -14275 5048
rect -14241 5014 -14207 5048
rect -14173 5014 -14139 5048
rect -14105 5014 -14071 5048
rect -14037 5014 -14003 5048
rect -13969 5014 -13935 5048
rect -13901 5014 -13867 5048
rect -13833 5014 -13799 5048
rect -13765 5014 -13731 5048
rect -13697 5014 -13663 5048
rect -13629 5014 -13595 5048
rect -13561 5014 -13527 5048
rect -13493 5014 -13459 5048
rect -13425 5014 -13391 5048
rect -13357 5014 -13323 5048
rect -13289 5014 -13255 5048
rect -13221 5014 -13187 5048
rect -13153 5014 -13119 5048
rect -13085 5014 -13051 5048
rect -13017 5014 -12983 5048
rect -12949 5014 -12915 5048
rect -12881 5014 -12847 5048
rect -12813 5014 -12779 5048
rect -12745 5014 -12711 5048
rect -12677 5014 -12643 5048
rect -12609 5014 -12575 5048
rect -12541 5014 -12507 5048
rect -12473 5014 -12439 5048
rect -12405 5014 -12371 5048
rect -12337 5014 -12303 5048
rect -12269 5014 -12235 5048
rect -12201 5014 -12167 5048
rect -12133 5014 -12099 5048
rect -12065 5014 -12031 5048
rect -11997 5014 -11963 5048
rect -11929 5014 -11895 5048
rect -11861 5014 -11827 5048
rect -11793 5014 -11759 5048
rect -11725 5014 -11691 5048
rect -11657 5014 -11623 5048
rect -11589 5014 -11555 5048
rect -11521 5014 -11487 5048
rect -11453 5014 -11419 5048
rect -11385 5014 -11351 5048
rect -11317 5014 -11283 5048
rect -11249 5014 -11215 5048
rect -11181 5014 -11147 5048
rect -11113 5014 -11079 5048
rect -11045 5014 -11011 5048
rect -10977 5014 -10943 5048
rect -10909 5014 -10875 5048
rect -10841 5014 -10807 5048
rect -10773 5014 -10739 5048
rect -10705 5014 -10671 5048
rect -10637 5014 -10603 5048
rect -10569 5014 -10535 5048
rect -10501 5014 -10467 5048
rect -10433 5014 -10399 5048
rect -10365 5014 -10331 5048
rect -10297 5014 -10263 5048
rect -10229 5014 -10195 5048
rect -10161 5014 -10127 5048
rect -10093 5014 -10059 5048
rect -10025 5014 -9991 5048
rect -9957 5014 -9923 5048
rect -9889 5014 -9855 5048
rect -9821 5014 -9787 5048
rect -9753 5014 -9719 5048
rect -9685 5014 -9651 5048
rect -9617 5014 -9583 5048
rect -9549 5014 -9515 5048
rect -9481 5014 -9447 5048
rect -9413 5014 -9379 5048
rect -9345 5014 -9311 5048
rect -9277 5014 -9243 5048
rect -9209 5014 -9175 5048
rect -9141 5014 -9107 5048
rect -9073 5014 -9039 5048
rect -9005 5014 -8971 5048
rect -8937 5014 -8903 5048
rect -8869 5014 -8835 5048
rect -8801 5014 -8767 5048
rect -8733 5014 -8699 5048
rect -8665 5014 -8631 5048
rect -8597 5014 -8563 5048
rect -8529 5014 -8495 5048
rect -8461 5014 -8427 5048
rect -8393 5014 -8359 5048
rect -8325 5014 -8291 5048
rect -8257 5014 -8223 5048
rect -8189 5014 -8155 5048
rect -8121 5014 -8087 5048
rect -8053 5014 -8019 5048
rect -7985 5014 -7951 5048
rect -7917 5014 -7883 5048
rect -7849 5014 -7815 5048
rect -7781 5014 -7747 5048
rect -7713 5014 -7679 5048
rect -7645 5014 -7611 5048
rect -7577 5014 -7543 5048
<< locali >>
rect -18121 8847 -18034 8881
rect -18000 8847 -17966 8881
rect -17932 8847 -17898 8881
rect -17864 8847 -17830 8881
rect -17796 8847 -17762 8881
rect -17728 8847 -17694 8881
rect -17660 8847 -17626 8881
rect -17592 8847 -17558 8881
rect -17524 8847 -17490 8881
rect -17456 8847 -17422 8881
rect -17388 8847 -17354 8881
rect -17320 8847 -17286 8881
rect -17252 8847 -17218 8881
rect -17184 8847 -17150 8881
rect -17116 8847 -17082 8881
rect -17048 8847 -17014 8881
rect -16980 8847 -16946 8881
rect -16912 8847 -16878 8881
rect -16844 8847 -16810 8881
rect -16776 8847 -16742 8881
rect -16708 8847 -16674 8881
rect -16640 8847 -16606 8881
rect -16572 8847 -16538 8881
rect -16504 8847 -16470 8881
rect -16436 8847 -16402 8881
rect -16368 8847 -16334 8881
rect -16300 8847 -16266 8881
rect -16232 8847 -16198 8881
rect -16164 8847 -16130 8881
rect -16096 8847 -16062 8881
rect -16028 8847 -15994 8881
rect -15960 8847 -15926 8881
rect -15892 8847 -15858 8881
rect -15824 8847 -15790 8881
rect -15756 8847 -15722 8881
rect -15688 8847 -15654 8881
rect -15620 8847 -15586 8881
rect -15552 8847 -15518 8881
rect -15484 8847 -15450 8881
rect -15416 8847 -15382 8881
rect -15348 8847 -15314 8881
rect -15280 8847 -15246 8881
rect -15212 8847 -15178 8881
rect -15144 8847 -15110 8881
rect -15076 8847 -15042 8881
rect -15008 8847 -14974 8881
rect -14940 8847 -14906 8881
rect -14872 8847 -14838 8881
rect -14804 8847 -14770 8881
rect -14736 8847 -14702 8881
rect -14668 8847 -14634 8881
rect -14600 8847 -14566 8881
rect -14532 8847 -14498 8881
rect -14464 8847 -14430 8881
rect -14396 8847 -14362 8881
rect -14328 8847 -14294 8881
rect -14260 8847 -14226 8881
rect -14192 8847 -14158 8881
rect -14124 8847 -14090 8881
rect -14056 8847 -14022 8881
rect -13988 8847 -13954 8881
rect -13920 8847 -13886 8881
rect -13852 8847 -13818 8881
rect -13784 8847 -13750 8881
rect -13716 8847 -13682 8881
rect -13648 8847 -13614 8881
rect -13580 8847 -13546 8881
rect -13512 8847 -13478 8881
rect -13444 8847 -13410 8881
rect -13376 8847 -13342 8881
rect -13308 8847 -13274 8881
rect -13240 8847 -13206 8881
rect -13172 8847 -13138 8881
rect -13104 8847 -13070 8881
rect -13036 8847 -13002 8881
rect -12968 8847 -12934 8881
rect -12900 8847 -12866 8881
rect -12832 8847 -12798 8881
rect -12764 8847 -12730 8881
rect -12696 8847 -12662 8881
rect -12628 8847 -12594 8881
rect -12560 8847 -12526 8881
rect -12492 8847 -12458 8881
rect -12424 8847 -12390 8881
rect -12356 8847 -12322 8881
rect -12288 8847 -12254 8881
rect -12220 8847 -12186 8881
rect -12152 8847 -12118 8881
rect -12084 8847 -12050 8881
rect -12016 8847 -11982 8881
rect -11948 8847 -11914 8881
rect -11880 8847 -11846 8881
rect -11812 8847 -11778 8881
rect -11744 8847 -11710 8881
rect -11676 8847 -11642 8881
rect -11608 8847 -11574 8881
rect -11540 8847 -11506 8881
rect -11472 8847 -11438 8881
rect -11404 8847 -11370 8881
rect -11336 8847 -11302 8881
rect -11268 8847 -11234 8881
rect -11200 8847 -11166 8881
rect -11132 8847 -11098 8881
rect -11064 8847 -11030 8881
rect -10996 8847 -10962 8881
rect -10928 8847 -10894 8881
rect -10860 8847 -10826 8881
rect -10792 8847 -10758 8881
rect -10724 8847 -10690 8881
rect -10656 8847 -10622 8881
rect -10588 8847 -10554 8881
rect -10520 8847 -10486 8881
rect -10452 8847 -10418 8881
rect -10384 8847 -10350 8881
rect -10316 8847 -10282 8881
rect -10248 8847 -10214 8881
rect -10180 8847 -10146 8881
rect -10112 8847 -10078 8881
rect -10044 8847 -10010 8881
rect -9976 8847 -9942 8881
rect -9908 8847 -9874 8881
rect -9840 8847 -9806 8881
rect -9772 8847 -9738 8881
rect -9704 8847 -9670 8881
rect -9636 8847 -9602 8881
rect -9568 8847 -9534 8881
rect -9500 8847 -9466 8881
rect -9432 8847 -9398 8881
rect -9364 8847 -9330 8881
rect -9296 8847 -9262 8881
rect -9228 8847 -9194 8881
rect -9160 8847 -9126 8881
rect -9092 8847 -9058 8881
rect -9024 8847 -8990 8881
rect -8956 8847 -8922 8881
rect -8888 8847 -8854 8881
rect -8820 8847 -8786 8881
rect -8752 8847 -8718 8881
rect -8684 8847 -8650 8881
rect -8616 8847 -8582 8881
rect -8548 8847 -8514 8881
rect -8480 8847 -8446 8881
rect -8412 8847 -8378 8881
rect -8344 8847 -8310 8881
rect -8276 8847 -8242 8881
rect -8208 8847 -8174 8881
rect -8140 8847 -8106 8881
rect -8072 8847 -8038 8881
rect -8004 8847 -7970 8881
rect -7936 8847 -7902 8881
rect -7868 8847 -7834 8881
rect -7800 8847 -7766 8881
rect -7732 8847 -7698 8881
rect -7664 8847 -7630 8881
rect -7596 8847 -7562 8881
rect -7528 8847 -7385 8881
rect -18121 8741 -18087 8847
rect -18121 8673 -18087 8707
rect -18121 8605 -18087 8639
rect -18121 8537 -18087 8571
rect -18121 8469 -18087 8503
rect -18121 8401 -18087 8435
rect -18121 8333 -18087 8367
rect -18121 8265 -18087 8299
rect -18121 8197 -18087 8231
rect -18121 8129 -18087 8163
rect -18121 8061 -18087 8095
rect -18121 7993 -18087 8027
rect -18121 7925 -18087 7959
rect -18121 7857 -18087 7891
rect -18121 7789 -18087 7823
rect -18121 7721 -18087 7755
rect -18121 7653 -18087 7687
rect -18121 7585 -18087 7619
rect -18121 7517 -18087 7551
rect -18121 7449 -18087 7483
rect -18121 7381 -18087 7415
rect -18121 7313 -18087 7347
rect -18121 7245 -18087 7279
rect -18121 7177 -18087 7211
rect -18121 7109 -18087 7143
rect -18121 7041 -18087 7075
rect -18121 6973 -18087 7007
rect -18121 6905 -18087 6939
rect -18121 6837 -18087 6871
rect -18121 6769 -18087 6803
rect -18121 6701 -18087 6735
rect -18121 6633 -18087 6667
rect -18121 6565 -18087 6599
rect -18121 6497 -18087 6531
rect -18121 6429 -18087 6463
rect -18121 6361 -18087 6395
rect -18121 6293 -18087 6327
rect -18121 6225 -18087 6259
rect -18121 6157 -18087 6191
rect -18121 6089 -18087 6123
rect -18121 6021 -18087 6055
rect -18121 5953 -18087 5987
rect -18121 5885 -18087 5919
rect -18121 5817 -18087 5851
rect -18121 5749 -18087 5783
rect -18121 5681 -18087 5715
rect -18121 5613 -18087 5647
rect -18121 5545 -18087 5579
rect -18121 5477 -18087 5511
rect -18121 5409 -18087 5443
rect -18121 5341 -18087 5375
rect -18121 5273 -18087 5307
rect -18121 5205 -18087 5239
rect -18121 5048 -18087 5171
rect -7419 8741 -7385 8847
rect -7419 8673 -7385 8707
rect -7419 8605 -7385 8639
rect -7419 8537 -7385 8571
rect -7419 8469 -7385 8503
rect -7419 8401 -7385 8435
rect -7419 8333 -7385 8367
rect -7419 8265 -7385 8299
rect -7419 8197 -7385 8231
rect -7419 8129 -7385 8163
rect -7419 8061 -7385 8095
rect -7419 7993 -7385 8027
rect -7419 7925 -7385 7959
rect -7419 7857 -7385 7891
rect -7419 7789 -7385 7823
rect -7419 7721 -7385 7755
rect -7419 7653 -7385 7687
rect -7419 7585 -7385 7619
rect -7419 7517 -7385 7551
rect -7419 7449 -7385 7483
rect -7419 7381 -7385 7415
rect -7419 7313 -7385 7347
rect -7419 7245 -7385 7279
rect -7419 7177 -7385 7211
rect -7419 7109 -7385 7143
rect -7419 7041 -7385 7075
rect -7419 6973 -7385 7007
rect -7419 6905 -7385 6939
rect -7419 6837 -7385 6871
rect -7419 6769 -7385 6803
rect -7419 6701 -7385 6735
rect -7419 6633 -7385 6667
rect -7419 6565 -7385 6599
rect -7419 6497 -7385 6531
rect -7419 6429 -7385 6463
rect -7419 6361 -7385 6395
rect -7419 6293 -7385 6327
rect -7419 6225 -7385 6259
rect -7419 6157 -7385 6191
rect -7419 6089 -7385 6123
rect -7419 6021 -7385 6055
rect -7419 5953 -7385 5987
rect -7419 5885 -7385 5919
rect -7419 5817 -7385 5851
rect -7419 5749 -7385 5783
rect -7419 5681 -7385 5715
rect -7419 5613 -7385 5647
rect -7419 5545 -7385 5579
rect -7419 5477 -7385 5511
rect -7419 5409 -7385 5443
rect -7419 5341 -7385 5375
rect -7419 5273 -7385 5307
rect -7419 5205 -7385 5239
rect -7419 5048 -7385 5171
rect -18121 5014 -17981 5048
rect -17947 5014 -17913 5048
rect -17879 5014 -17845 5048
rect -17811 5014 -17777 5048
rect -17743 5014 -17709 5048
rect -17675 5014 -17641 5048
rect -17607 5014 -17573 5048
rect -17539 5014 -17505 5048
rect -17471 5014 -17437 5048
rect -17403 5014 -17369 5048
rect -17335 5014 -17301 5048
rect -17267 5014 -17233 5048
rect -17199 5014 -17165 5048
rect -17131 5014 -17097 5048
rect -17063 5014 -17029 5048
rect -16995 5014 -16961 5048
rect -16927 5014 -16893 5048
rect -16859 5014 -16825 5048
rect -16791 5014 -16757 5048
rect -16723 5014 -16689 5048
rect -16655 5014 -16621 5048
rect -16587 5014 -16553 5048
rect -16519 5014 -16485 5048
rect -16451 5014 -16417 5048
rect -16383 5014 -16349 5048
rect -16315 5014 -16281 5048
rect -16247 5014 -16213 5048
rect -16179 5014 -16145 5048
rect -16111 5014 -16077 5048
rect -16043 5014 -16009 5048
rect -15975 5014 -15941 5048
rect -15907 5014 -15873 5048
rect -15839 5014 -15805 5048
rect -15771 5014 -15737 5048
rect -15703 5014 -15669 5048
rect -15635 5014 -15601 5048
rect -15567 5014 -15533 5048
rect -15499 5014 -15465 5048
rect -15431 5014 -15397 5048
rect -15363 5014 -15329 5048
rect -15295 5014 -15261 5048
rect -15227 5014 -15193 5048
rect -15159 5014 -15125 5048
rect -15091 5014 -15057 5048
rect -15023 5014 -14989 5048
rect -14955 5014 -14921 5048
rect -14887 5014 -14853 5048
rect -14819 5014 -14785 5048
rect -14751 5014 -14717 5048
rect -14683 5014 -14649 5048
rect -14615 5014 -14581 5048
rect -14547 5014 -14513 5048
rect -14479 5014 -14445 5048
rect -14411 5014 -14377 5048
rect -14343 5014 -14309 5048
rect -14275 5014 -14241 5048
rect -14207 5014 -14173 5048
rect -14139 5014 -14105 5048
rect -14071 5014 -14037 5048
rect -14003 5014 -13969 5048
rect -13935 5014 -13901 5048
rect -13867 5014 -13833 5048
rect -13799 5014 -13765 5048
rect -13731 5014 -13697 5048
rect -13663 5014 -13629 5048
rect -13595 5014 -13561 5048
rect -13527 5014 -13493 5048
rect -13459 5014 -13425 5048
rect -13391 5014 -13357 5048
rect -13323 5014 -13289 5048
rect -13255 5014 -13221 5048
rect -13187 5014 -13153 5048
rect -13119 5014 -13085 5048
rect -13051 5014 -13017 5048
rect -12983 5014 -12949 5048
rect -12915 5014 -12881 5048
rect -12847 5014 -12813 5048
rect -12779 5014 -12745 5048
rect -12711 5014 -12677 5048
rect -12643 5014 -12609 5048
rect -12575 5014 -12541 5048
rect -12507 5014 -12473 5048
rect -12439 5014 -12405 5048
rect -12371 5014 -12337 5048
rect -12303 5014 -12269 5048
rect -12235 5014 -12201 5048
rect -12167 5014 -12133 5048
rect -12099 5014 -12065 5048
rect -12031 5014 -11997 5048
rect -11963 5014 -11929 5048
rect -11895 5014 -11861 5048
rect -11827 5014 -11793 5048
rect -11759 5014 -11725 5048
rect -11691 5014 -11657 5048
rect -11623 5014 -11589 5048
rect -11555 5014 -11521 5048
rect -11487 5014 -11453 5048
rect -11419 5014 -11385 5048
rect -11351 5014 -11317 5048
rect -11283 5014 -11249 5048
rect -11215 5014 -11181 5048
rect -11147 5014 -11113 5048
rect -11079 5014 -11045 5048
rect -11011 5014 -10977 5048
rect -10943 5014 -10909 5048
rect -10875 5014 -10841 5048
rect -10807 5014 -10773 5048
rect -10739 5014 -10705 5048
rect -10671 5014 -10637 5048
rect -10603 5014 -10569 5048
rect -10535 5014 -10501 5048
rect -10467 5014 -10433 5048
rect -10399 5014 -10365 5048
rect -10331 5014 -10297 5048
rect -10263 5014 -10229 5048
rect -10195 5014 -10161 5048
rect -10127 5014 -10093 5048
rect -10059 5014 -10025 5048
rect -9991 5014 -9957 5048
rect -9923 5014 -9889 5048
rect -9855 5014 -9821 5048
rect -9787 5014 -9753 5048
rect -9719 5014 -9685 5048
rect -9651 5014 -9617 5048
rect -9583 5014 -9549 5048
rect -9515 5014 -9481 5048
rect -9447 5014 -9413 5048
rect -9379 5014 -9345 5048
rect -9311 5014 -9277 5048
rect -9243 5014 -9209 5048
rect -9175 5014 -9141 5048
rect -9107 5014 -9073 5048
rect -9039 5014 -9005 5048
rect -8971 5014 -8937 5048
rect -8903 5014 -8869 5048
rect -8835 5014 -8801 5048
rect -8767 5014 -8733 5048
rect -8699 5014 -8665 5048
rect -8631 5014 -8597 5048
rect -8563 5014 -8529 5048
rect -8495 5014 -8461 5048
rect -8427 5014 -8393 5048
rect -8359 5014 -8325 5048
rect -8291 5014 -8257 5048
rect -8223 5014 -8189 5048
rect -8155 5014 -8121 5048
rect -8087 5014 -8053 5048
rect -8019 5014 -7985 5048
rect -7951 5014 -7917 5048
rect -7883 5014 -7849 5048
rect -7815 5014 -7781 5048
rect -7747 5014 -7713 5048
rect -7679 5014 -7645 5048
rect -7611 5014 -7577 5048
rect -7543 5014 -7385 5048
<< properties >>
string path -90.785 44.320 -37.010 44.320 -37.010 25.155 -90.520 25.155 -90.520 44.320 
<< end >>
