magic
tech sky130A
magscale 1 2
timestamp 1715625863
<< nwell >>
rect -425 -284 425 284
<< pmos >>
rect -229 -136 -29 64
rect 29 -136 229 64
<< pdiff >>
rect -287 49 -229 64
rect -287 15 -275 49
rect -241 15 -229 49
rect -287 -19 -229 15
rect -287 -53 -275 -19
rect -241 -53 -229 -19
rect -287 -87 -229 -53
rect -287 -121 -275 -87
rect -241 -121 -229 -87
rect -287 -136 -229 -121
rect -29 49 29 64
rect -29 15 -17 49
rect 17 15 29 49
rect -29 -19 29 15
rect -29 -53 -17 -19
rect 17 -53 29 -19
rect -29 -87 29 -53
rect -29 -121 -17 -87
rect 17 -121 29 -87
rect -29 -136 29 -121
rect 229 49 287 64
rect 229 15 241 49
rect 275 15 287 49
rect 229 -19 287 15
rect 229 -53 241 -19
rect 275 -53 287 -19
rect 229 -87 287 -53
rect 229 -121 241 -87
rect 275 -121 287 -87
rect 229 -136 287 -121
<< pdiffc >>
rect -275 15 -241 49
rect -275 -53 -241 -19
rect -275 -121 -241 -87
rect -17 15 17 49
rect -17 -53 17 -19
rect -17 -121 17 -87
rect 241 15 275 49
rect 241 -53 275 -19
rect 241 -121 275 -87
<< nsubdiff >>
rect -389 214 -289 248
rect -255 214 -221 248
rect -187 214 -153 248
rect -119 214 -85 248
rect -51 214 -17 248
rect 17 214 51 248
rect 85 214 119 248
rect 153 214 187 248
rect 221 214 255 248
rect 289 214 389 248
rect -389 119 -355 214
rect -389 51 -355 85
rect 355 119 389 214
rect -389 -17 -355 17
rect -389 -85 -355 -51
rect -389 -214 -355 -119
rect 355 51 389 85
rect 355 -17 389 17
rect 355 -85 389 -51
rect 355 -214 389 -119
rect -389 -248 -289 -214
rect -255 -248 -221 -214
rect -187 -248 -153 -214
rect -119 -248 -85 -214
rect -51 -248 -17 -214
rect 17 -248 51 -214
rect 85 -248 119 -214
rect 153 -248 187 -214
rect 221 -248 255 -214
rect 289 -248 389 -214
<< nsubdiffcont >>
rect -289 214 -255 248
rect -221 214 -187 248
rect -153 214 -119 248
rect -85 214 -51 248
rect -17 214 17 248
rect 51 214 85 248
rect 119 214 153 248
rect 187 214 221 248
rect 255 214 289 248
rect -389 85 -355 119
rect 355 85 389 119
rect -389 17 -355 51
rect -389 -51 -355 -17
rect -389 -119 -355 -85
rect 355 17 389 51
rect 355 -51 389 -17
rect 355 -119 389 -85
rect -289 -248 -255 -214
rect -221 -248 -187 -214
rect -153 -248 -119 -214
rect -85 -248 -51 -214
rect -17 -248 17 -214
rect 51 -248 85 -214
rect 119 -248 153 -214
rect 187 -248 221 -214
rect 255 -248 289 -214
<< poly >>
rect -229 145 -29 161
rect -229 111 -180 145
rect -146 111 -112 145
rect -78 111 -29 145
rect -229 64 -29 111
rect 29 145 229 161
rect 29 111 78 145
rect 112 111 146 145
rect 180 111 229 145
rect 29 64 229 111
rect -229 -162 -29 -136
rect 29 -162 229 -136
<< polycont >>
rect -180 111 -146 145
rect -112 111 -78 145
rect 78 111 112 145
rect 146 111 180 145
<< locali >>
rect -389 214 -289 248
rect -255 214 -221 248
rect -187 214 -153 248
rect -119 214 -85 248
rect -51 214 -17 248
rect 17 214 51 248
rect 85 214 119 248
rect 153 214 187 248
rect 221 214 255 248
rect 289 214 389 248
rect -389 119 -355 214
rect -229 111 -182 145
rect -146 111 -112 145
rect -76 111 -29 145
rect 29 111 76 145
rect 112 111 146 145
rect 182 111 229 145
rect 355 119 389 214
rect -389 51 -355 85
rect -389 -17 -355 17
rect -389 -85 -355 -51
rect -389 -214 -355 -119
rect -275 49 -241 68
rect -275 -19 -241 -17
rect -275 -55 -241 -53
rect -275 -140 -241 -121
rect -17 49 17 68
rect -17 -19 17 -17
rect -17 -55 17 -53
rect -17 -140 17 -121
rect 241 49 275 68
rect 241 -19 275 -17
rect 241 -55 275 -53
rect 241 -140 275 -121
rect 355 51 389 85
rect 355 -17 389 17
rect 355 -85 389 -51
rect 355 -214 389 -119
rect -389 -248 -289 -214
rect -255 -248 -221 -214
rect -187 -248 -153 -214
rect -119 -248 -85 -214
rect -51 -248 -17 -214
rect 17 -248 51 -214
rect 85 -248 119 -214
rect 153 -248 187 -214
rect 221 -248 255 -214
rect 289 -248 389 -214
<< viali >>
rect -182 111 -180 145
rect -180 111 -148 145
rect -110 111 -78 145
rect -78 111 -76 145
rect 76 111 78 145
rect 78 111 110 145
rect 148 111 180 145
rect 180 111 182 145
rect -275 15 -241 17
rect -275 -17 -241 15
rect -275 -87 -241 -55
rect -275 -89 -241 -87
rect -17 15 17 17
rect -17 -17 17 15
rect -17 -87 17 -55
rect -17 -89 17 -87
rect 241 15 275 17
rect 241 -17 275 15
rect 241 -87 275 -55
rect 241 -89 275 -87
<< metal1 >>
rect -225 145 -33 151
rect -225 111 -182 145
rect -148 111 -110 145
rect -76 111 -33 145
rect -225 105 -33 111
rect 33 145 225 151
rect 33 111 76 145
rect 110 111 148 145
rect 182 111 225 145
rect 33 105 225 111
rect -281 17 -235 64
rect -281 -17 -275 17
rect -241 -17 -235 17
rect -281 -55 -235 -17
rect -281 -89 -275 -55
rect -241 -89 -235 -55
rect -281 -136 -235 -89
rect -23 17 23 64
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -136 23 -89
rect 235 17 281 64
rect 235 -17 241 17
rect 275 -17 281 17
rect 235 -55 281 -17
rect 235 -89 241 -55
rect 275 -89 281 -55
rect 235 -136 281 -89
<< properties >>
string FIXED_BBOX -372 -231 372 231
<< end >>
