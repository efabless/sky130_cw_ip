magic
tech sky130A
magscale 1 2
timestamp 1715010268
<< nwell >>
rect -194 -148 194 114
<< pmoslvt >>
rect -100 -86 100 14
<< pdiff >>
rect -158 -19 -100 14
rect -158 -53 -146 -19
rect -112 -53 -100 -19
rect -158 -86 -100 -53
rect 100 -19 158 14
rect 100 -53 112 -19
rect 146 -53 158 -19
rect 100 -86 158 -53
<< pdiffc >>
rect -146 -53 -112 -19
rect 112 -53 146 -19
<< poly >>
rect -100 95 100 111
rect -100 61 -51 95
rect -17 61 17 95
rect 51 61 100 95
rect -100 14 100 61
rect -100 -112 100 -86
<< polycont >>
rect -51 61 -17 95
rect 17 61 51 95
<< locali >>
rect -100 61 -53 95
rect -17 61 17 95
rect 53 61 100 95
rect -146 -19 -112 18
rect -146 -90 -112 -53
rect 112 -19 146 18
rect 112 -90 146 -53
<< viali >>
rect -53 61 -51 95
rect -51 61 -19 95
rect 19 61 51 95
rect 51 61 53 95
rect -146 -53 -112 -19
rect 112 -53 146 -19
<< metal1 >>
rect -96 95 96 101
rect -96 61 -53 95
rect -19 61 19 95
rect 53 61 96 95
rect -96 55 96 61
rect -152 -19 -106 14
rect -152 -53 -146 -19
rect -112 -53 -106 -19
rect -152 -86 -106 -53
rect 106 -19 152 14
rect 106 -53 112 -19
rect 146 -53 152 -19
rect 106 -86 152 -53
<< end >>
