magic
tech sky130A
magscale 1 2
timestamp 1715010268
<< pwell >>
rect -415 -269 415 269
<< nmos >>
rect -229 -131 -29 69
rect 29 -131 229 69
<< ndiff >>
rect -287 54 -229 69
rect -287 20 -275 54
rect -241 20 -229 54
rect -287 -14 -229 20
rect -287 -48 -275 -14
rect -241 -48 -229 -14
rect -287 -82 -229 -48
rect -287 -116 -275 -82
rect -241 -116 -229 -82
rect -287 -131 -229 -116
rect -29 54 29 69
rect -29 20 -17 54
rect 17 20 29 54
rect -29 -14 29 20
rect -29 -48 -17 -14
rect 17 -48 29 -14
rect -29 -82 29 -48
rect -29 -116 -17 -82
rect 17 -116 29 -82
rect -29 -131 29 -116
rect 229 54 287 69
rect 229 20 241 54
rect 275 20 287 54
rect 229 -14 287 20
rect 229 -48 241 -14
rect 275 -48 287 -14
rect 229 -82 287 -48
rect 229 -116 241 -82
rect 275 -116 287 -82
rect 229 -131 287 -116
<< ndiffc >>
rect -275 20 -241 54
rect -275 -48 -241 -14
rect -275 -116 -241 -82
rect -17 20 17 54
rect -17 -48 17 -14
rect -17 -116 17 -82
rect 241 20 275 54
rect 241 -48 275 -14
rect 241 -116 275 -82
<< psubdiff >>
rect -389 209 -289 243
rect -255 209 -221 243
rect -187 209 -153 243
rect -119 209 -85 243
rect -51 209 -17 243
rect 17 209 51 243
rect 85 209 119 243
rect 153 209 187 243
rect 221 209 255 243
rect 289 209 389 243
rect -389 119 -355 209
rect -389 51 -355 85
rect 355 119 389 209
rect -389 -17 -355 17
rect -389 -85 -355 -51
rect -389 -209 -355 -119
rect 355 51 389 85
rect 355 -17 389 17
rect 355 -85 389 -51
rect 355 -209 389 -119
rect -389 -243 -289 -209
rect -255 -243 -221 -209
rect -187 -243 -153 -209
rect -119 -243 -85 -209
rect -51 -243 -17 -209
rect 17 -243 51 -209
rect 85 -243 119 -209
rect 153 -243 187 -209
rect 221 -243 255 -209
rect 289 -243 389 -209
<< psubdiffcont >>
rect -289 209 -255 243
rect -221 209 -187 243
rect -153 209 -119 243
rect -85 209 -51 243
rect -17 209 17 243
rect 51 209 85 243
rect 119 209 153 243
rect 187 209 221 243
rect 255 209 289 243
rect -389 85 -355 119
rect 355 85 389 119
rect -389 17 -355 51
rect -389 -51 -355 -17
rect -389 -119 -355 -85
rect 355 17 389 51
rect 355 -51 389 -17
rect 355 -119 389 -85
rect -289 -243 -255 -209
rect -221 -243 -187 -209
rect -153 -243 -119 -209
rect -85 -243 -51 -209
rect -17 -243 17 -209
rect 51 -243 85 -209
rect 119 -243 153 -209
rect 187 -243 221 -209
rect 255 -243 289 -209
<< poly >>
rect -229 141 -29 157
rect -229 107 -180 141
rect -146 107 -112 141
rect -78 107 -29 141
rect -229 69 -29 107
rect 29 141 229 157
rect 29 107 78 141
rect 112 107 146 141
rect 180 107 229 141
rect 29 69 229 107
rect -229 -157 -29 -131
rect 29 -157 229 -131
<< polycont >>
rect -180 107 -146 141
rect -112 107 -78 141
rect 78 107 112 141
rect 146 107 180 141
<< locali >>
rect -389 209 -289 243
rect -255 209 -221 243
rect -187 209 -153 243
rect -119 209 -85 243
rect -51 209 -17 243
rect 17 209 51 243
rect 85 209 119 243
rect 153 209 187 243
rect 221 209 255 243
rect 289 209 389 243
rect -389 119 -355 209
rect -229 107 -182 141
rect -146 107 -112 141
rect -76 107 -29 141
rect 29 107 76 141
rect 112 107 146 141
rect 182 107 229 141
rect 355 119 389 209
rect -389 51 -355 85
rect -389 -17 -355 17
rect -389 -85 -355 -51
rect -389 -209 -355 -119
rect -275 54 -241 73
rect -275 -14 -241 -12
rect -275 -50 -241 -48
rect -275 -135 -241 -116
rect -17 54 17 73
rect -17 -14 17 -12
rect -17 -50 17 -48
rect -17 -135 17 -116
rect 241 54 275 73
rect 241 -14 275 -12
rect 241 -50 275 -48
rect 241 -135 275 -116
rect 355 51 389 85
rect 355 -17 389 17
rect 355 -85 389 -51
rect 355 -209 389 -119
rect -389 -243 -289 -209
rect -255 -243 -221 -209
rect -187 -243 -153 -209
rect -119 -243 -85 -209
rect -51 -243 -17 -209
rect 17 -243 51 -209
rect 85 -243 119 -209
rect 153 -243 187 -209
rect 221 -243 255 -209
rect 289 -243 389 -209
<< viali >>
rect -182 107 -180 141
rect -180 107 -148 141
rect -110 107 -78 141
rect -78 107 -76 141
rect 76 107 78 141
rect 78 107 110 141
rect 148 107 180 141
rect 180 107 182 141
rect -275 20 -241 22
rect -275 -12 -241 20
rect -275 -82 -241 -50
rect -275 -84 -241 -82
rect -17 20 17 22
rect -17 -12 17 20
rect -17 -82 17 -50
rect -17 -84 17 -82
rect 241 20 275 22
rect 241 -12 275 20
rect 241 -82 275 -50
rect 241 -84 275 -82
<< metal1 >>
rect -225 141 -33 147
rect -225 107 -182 141
rect -148 107 -110 141
rect -76 107 -33 141
rect -225 101 -33 107
rect 33 141 225 147
rect 33 107 76 141
rect 110 107 148 141
rect 182 107 225 141
rect 33 101 225 107
rect -281 22 -235 69
rect -281 -12 -275 22
rect -241 -12 -235 22
rect -281 -50 -235 -12
rect -281 -84 -275 -50
rect -241 -84 -235 -50
rect -281 -131 -235 -84
rect -23 22 23 69
rect -23 -12 -17 22
rect 17 -12 23 22
rect -23 -50 23 -12
rect -23 -84 -17 -50
rect 17 -84 23 -50
rect -23 -131 23 -84
rect 235 22 281 69
rect 235 -12 241 22
rect 275 -12 281 22
rect 235 -50 281 -12
rect 235 -84 241 -50
rect 275 -84 281 -50
rect 235 -131 281 -84
<< properties >>
string FIXED_BBOX -372 -226 372 226
<< end >>
