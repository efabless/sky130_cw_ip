magic
tech sky130A
magscale 1 2
timestamp 1715625863
<< pwell >>
rect -14705 5391 -9167 5477
rect -14705 2733 -14619 5391
rect -9253 2733 -9167 5391
rect -14705 2647 -9167 2733
<< psubdiff >>
rect -14679 5417 -14521 5451
rect -14487 5417 -14453 5451
rect -14419 5417 -14385 5451
rect -14351 5417 -14317 5451
rect -14283 5417 -14249 5451
rect -14215 5417 -14181 5451
rect -14147 5417 -14113 5451
rect -14079 5417 -14045 5451
rect -14011 5417 -13977 5451
rect -13943 5417 -13909 5451
rect -13875 5417 -13841 5451
rect -13807 5417 -13773 5451
rect -13739 5417 -13705 5451
rect -13671 5417 -13637 5451
rect -13603 5417 -13569 5451
rect -13535 5417 -13501 5451
rect -13467 5417 -13433 5451
rect -13399 5417 -13365 5451
rect -13331 5417 -13297 5451
rect -13263 5417 -13229 5451
rect -13195 5417 -13161 5451
rect -13127 5417 -13093 5451
rect -13059 5417 -13025 5451
rect -12991 5417 -12957 5451
rect -12923 5417 -12889 5451
rect -12855 5417 -12821 5451
rect -12787 5417 -12753 5451
rect -12719 5417 -12685 5451
rect -12651 5417 -12617 5451
rect -12583 5417 -12549 5451
rect -12515 5417 -12481 5451
rect -12447 5417 -12413 5451
rect -12379 5417 -12345 5451
rect -12311 5417 -12277 5451
rect -12243 5417 -12209 5451
rect -12175 5417 -12141 5451
rect -12107 5417 -12073 5451
rect -12039 5417 -12005 5451
rect -11971 5417 -11937 5451
rect -11903 5417 -11869 5451
rect -11835 5417 -11801 5451
rect -11767 5417 -11733 5451
rect -11699 5417 -11665 5451
rect -11631 5417 -11597 5451
rect -11563 5417 -11529 5451
rect -11495 5417 -11461 5451
rect -11427 5417 -11393 5451
rect -11359 5417 -11325 5451
rect -11291 5417 -11257 5451
rect -11223 5417 -11189 5451
rect -11155 5417 -11121 5451
rect -11087 5417 -11053 5451
rect -11019 5417 -10985 5451
rect -10951 5417 -10917 5451
rect -10883 5417 -10849 5451
rect -10815 5417 -10781 5451
rect -10747 5417 -10713 5451
rect -10679 5417 -10645 5451
rect -10611 5417 -10577 5451
rect -10543 5417 -10509 5451
rect -10475 5417 -10441 5451
rect -10407 5417 -10373 5451
rect -10339 5417 -10305 5451
rect -10271 5417 -10237 5451
rect -10203 5417 -10169 5451
rect -10135 5417 -10101 5451
rect -10067 5417 -10033 5451
rect -9999 5417 -9965 5451
rect -9931 5417 -9897 5451
rect -9863 5417 -9829 5451
rect -9795 5417 -9761 5451
rect -9727 5417 -9693 5451
rect -9659 5417 -9625 5451
rect -9591 5417 -9557 5451
rect -9523 5417 -9489 5451
rect -9455 5417 -9193 5451
rect -14679 5251 -14645 5417
rect -14679 5183 -14645 5217
rect -14679 5115 -14645 5149
rect -14679 5047 -14645 5081
rect -14679 4979 -14645 5013
rect -14679 4911 -14645 4945
rect -14679 4843 -14645 4877
rect -14679 4775 -14645 4809
rect -14679 4707 -14645 4741
rect -14679 4639 -14645 4673
rect -14679 4571 -14645 4605
rect -14679 4503 -14645 4537
rect -14679 4435 -14645 4469
rect -14679 4367 -14645 4401
rect -14679 4299 -14645 4333
rect -14679 4231 -14645 4265
rect -14679 4163 -14645 4197
rect -14679 4095 -14645 4129
rect -14679 4027 -14645 4061
rect -14679 3959 -14645 3993
rect -14679 3891 -14645 3925
rect -14679 3823 -14645 3857
rect -14679 3755 -14645 3789
rect -14679 3687 -14645 3721
rect -14679 3619 -14645 3653
rect -14679 3551 -14645 3585
rect -14679 3483 -14645 3517
rect -14679 3415 -14645 3449
rect -14679 3347 -14645 3381
rect -14679 3279 -14645 3313
rect -14679 3211 -14645 3245
rect -14679 3143 -14645 3177
rect -14679 3075 -14645 3109
rect -14679 3007 -14645 3041
rect -14679 2939 -14645 2973
rect -14679 2707 -14645 2905
rect -9227 5251 -9193 5417
rect -9227 5183 -9193 5217
rect -9227 5115 -9193 5149
rect -9227 5047 -9193 5081
rect -9227 4979 -9193 5013
rect -9227 4911 -9193 4945
rect -9227 4843 -9193 4877
rect -9227 4775 -9193 4809
rect -9227 4707 -9193 4741
rect -9227 4639 -9193 4673
rect -9227 4571 -9193 4605
rect -9227 4503 -9193 4537
rect -9227 4435 -9193 4469
rect -9227 4367 -9193 4401
rect -9227 4299 -9193 4333
rect -9227 4231 -9193 4265
rect -9227 4163 -9193 4197
rect -9227 4095 -9193 4129
rect -9227 4027 -9193 4061
rect -9227 3959 -9193 3993
rect -9227 3891 -9193 3925
rect -9227 3823 -9193 3857
rect -9227 3755 -9193 3789
rect -9227 3687 -9193 3721
rect -9227 3619 -9193 3653
rect -9227 3551 -9193 3585
rect -9227 3483 -9193 3517
rect -9227 3415 -9193 3449
rect -9227 3347 -9193 3381
rect -9227 3279 -9193 3313
rect -9227 3211 -9193 3245
rect -9227 3143 -9193 3177
rect -9227 3075 -9193 3109
rect -9227 3007 -9193 3041
rect -9227 2939 -9193 2973
rect -9227 2707 -9193 2905
rect -14679 2673 -14479 2707
rect -14445 2673 -14411 2707
rect -14377 2673 -14343 2707
rect -14309 2673 -14275 2707
rect -14241 2673 -14207 2707
rect -14173 2673 -14139 2707
rect -14105 2673 -14071 2707
rect -14037 2673 -14003 2707
rect -13969 2673 -13935 2707
rect -13901 2673 -13867 2707
rect -13833 2673 -13799 2707
rect -13765 2673 -13731 2707
rect -13697 2673 -13663 2707
rect -13629 2673 -13595 2707
rect -13561 2673 -13527 2707
rect -13493 2673 -13459 2707
rect -13425 2673 -13391 2707
rect -13357 2673 -13323 2707
rect -13289 2673 -13255 2707
rect -13221 2673 -13187 2707
rect -13153 2673 -13119 2707
rect -13085 2673 -13051 2707
rect -13017 2673 -12983 2707
rect -12949 2673 -12915 2707
rect -12881 2673 -12847 2707
rect -12813 2673 -12779 2707
rect -12745 2673 -12711 2707
rect -12677 2673 -12643 2707
rect -12609 2673 -12575 2707
rect -12541 2673 -12507 2707
rect -12473 2673 -12439 2707
rect -12405 2673 -12371 2707
rect -12337 2673 -12303 2707
rect -12269 2673 -12235 2707
rect -12201 2673 -12167 2707
rect -12133 2673 -12099 2707
rect -12065 2673 -12031 2707
rect -11997 2673 -11963 2707
rect -11929 2673 -11895 2707
rect -11861 2673 -11827 2707
rect -11793 2673 -11759 2707
rect -11725 2673 -11691 2707
rect -11657 2673 -11623 2707
rect -11589 2673 -11555 2707
rect -11521 2673 -11487 2707
rect -11453 2673 -11419 2707
rect -11385 2673 -11351 2707
rect -11317 2673 -11283 2707
rect -11249 2673 -11215 2707
rect -11181 2673 -11147 2707
rect -11113 2673 -11079 2707
rect -11045 2673 -11011 2707
rect -10977 2673 -10943 2707
rect -10909 2673 -10875 2707
rect -10841 2673 -10807 2707
rect -10773 2673 -10739 2707
rect -10705 2673 -10671 2707
rect -10637 2673 -10603 2707
rect -10569 2673 -10535 2707
rect -10501 2673 -10467 2707
rect -10433 2673 -10399 2707
rect -10365 2673 -10331 2707
rect -10297 2673 -10263 2707
rect -10229 2673 -10195 2707
rect -10161 2673 -10127 2707
rect -10093 2673 -10059 2707
rect -10025 2673 -9991 2707
rect -9957 2673 -9923 2707
rect -9889 2673 -9855 2707
rect -9821 2673 -9787 2707
rect -9753 2673 -9719 2707
rect -9685 2673 -9651 2707
rect -9617 2673 -9583 2707
rect -9549 2673 -9515 2707
rect -9481 2673 -9447 2707
rect -9413 2673 -9193 2707
<< psubdiffcont >>
rect -14521 5417 -14487 5451
rect -14453 5417 -14419 5451
rect -14385 5417 -14351 5451
rect -14317 5417 -14283 5451
rect -14249 5417 -14215 5451
rect -14181 5417 -14147 5451
rect -14113 5417 -14079 5451
rect -14045 5417 -14011 5451
rect -13977 5417 -13943 5451
rect -13909 5417 -13875 5451
rect -13841 5417 -13807 5451
rect -13773 5417 -13739 5451
rect -13705 5417 -13671 5451
rect -13637 5417 -13603 5451
rect -13569 5417 -13535 5451
rect -13501 5417 -13467 5451
rect -13433 5417 -13399 5451
rect -13365 5417 -13331 5451
rect -13297 5417 -13263 5451
rect -13229 5417 -13195 5451
rect -13161 5417 -13127 5451
rect -13093 5417 -13059 5451
rect -13025 5417 -12991 5451
rect -12957 5417 -12923 5451
rect -12889 5417 -12855 5451
rect -12821 5417 -12787 5451
rect -12753 5417 -12719 5451
rect -12685 5417 -12651 5451
rect -12617 5417 -12583 5451
rect -12549 5417 -12515 5451
rect -12481 5417 -12447 5451
rect -12413 5417 -12379 5451
rect -12345 5417 -12311 5451
rect -12277 5417 -12243 5451
rect -12209 5417 -12175 5451
rect -12141 5417 -12107 5451
rect -12073 5417 -12039 5451
rect -12005 5417 -11971 5451
rect -11937 5417 -11903 5451
rect -11869 5417 -11835 5451
rect -11801 5417 -11767 5451
rect -11733 5417 -11699 5451
rect -11665 5417 -11631 5451
rect -11597 5417 -11563 5451
rect -11529 5417 -11495 5451
rect -11461 5417 -11427 5451
rect -11393 5417 -11359 5451
rect -11325 5417 -11291 5451
rect -11257 5417 -11223 5451
rect -11189 5417 -11155 5451
rect -11121 5417 -11087 5451
rect -11053 5417 -11019 5451
rect -10985 5417 -10951 5451
rect -10917 5417 -10883 5451
rect -10849 5417 -10815 5451
rect -10781 5417 -10747 5451
rect -10713 5417 -10679 5451
rect -10645 5417 -10611 5451
rect -10577 5417 -10543 5451
rect -10509 5417 -10475 5451
rect -10441 5417 -10407 5451
rect -10373 5417 -10339 5451
rect -10305 5417 -10271 5451
rect -10237 5417 -10203 5451
rect -10169 5417 -10135 5451
rect -10101 5417 -10067 5451
rect -10033 5417 -9999 5451
rect -9965 5417 -9931 5451
rect -9897 5417 -9863 5451
rect -9829 5417 -9795 5451
rect -9761 5417 -9727 5451
rect -9693 5417 -9659 5451
rect -9625 5417 -9591 5451
rect -9557 5417 -9523 5451
rect -9489 5417 -9455 5451
rect -14679 5217 -14645 5251
rect -14679 5149 -14645 5183
rect -14679 5081 -14645 5115
rect -14679 5013 -14645 5047
rect -14679 4945 -14645 4979
rect -14679 4877 -14645 4911
rect -14679 4809 -14645 4843
rect -14679 4741 -14645 4775
rect -14679 4673 -14645 4707
rect -14679 4605 -14645 4639
rect -14679 4537 -14645 4571
rect -14679 4469 -14645 4503
rect -14679 4401 -14645 4435
rect -14679 4333 -14645 4367
rect -14679 4265 -14645 4299
rect -14679 4197 -14645 4231
rect -14679 4129 -14645 4163
rect -14679 4061 -14645 4095
rect -14679 3993 -14645 4027
rect -14679 3925 -14645 3959
rect -14679 3857 -14645 3891
rect -14679 3789 -14645 3823
rect -14679 3721 -14645 3755
rect -14679 3653 -14645 3687
rect -14679 3585 -14645 3619
rect -14679 3517 -14645 3551
rect -14679 3449 -14645 3483
rect -14679 3381 -14645 3415
rect -14679 3313 -14645 3347
rect -14679 3245 -14645 3279
rect -14679 3177 -14645 3211
rect -14679 3109 -14645 3143
rect -14679 3041 -14645 3075
rect -14679 2973 -14645 3007
rect -14679 2905 -14645 2939
rect -9227 5217 -9193 5251
rect -9227 5149 -9193 5183
rect -9227 5081 -9193 5115
rect -9227 5013 -9193 5047
rect -9227 4945 -9193 4979
rect -9227 4877 -9193 4911
rect -9227 4809 -9193 4843
rect -9227 4741 -9193 4775
rect -9227 4673 -9193 4707
rect -9227 4605 -9193 4639
rect -9227 4537 -9193 4571
rect -9227 4469 -9193 4503
rect -9227 4401 -9193 4435
rect -9227 4333 -9193 4367
rect -9227 4265 -9193 4299
rect -9227 4197 -9193 4231
rect -9227 4129 -9193 4163
rect -9227 4061 -9193 4095
rect -9227 3993 -9193 4027
rect -9227 3925 -9193 3959
rect -9227 3857 -9193 3891
rect -9227 3789 -9193 3823
rect -9227 3721 -9193 3755
rect -9227 3653 -9193 3687
rect -9227 3585 -9193 3619
rect -9227 3517 -9193 3551
rect -9227 3449 -9193 3483
rect -9227 3381 -9193 3415
rect -9227 3313 -9193 3347
rect -9227 3245 -9193 3279
rect -9227 3177 -9193 3211
rect -9227 3109 -9193 3143
rect -9227 3041 -9193 3075
rect -9227 2973 -9193 3007
rect -9227 2905 -9193 2939
rect -14479 2673 -14445 2707
rect -14411 2673 -14377 2707
rect -14343 2673 -14309 2707
rect -14275 2673 -14241 2707
rect -14207 2673 -14173 2707
rect -14139 2673 -14105 2707
rect -14071 2673 -14037 2707
rect -14003 2673 -13969 2707
rect -13935 2673 -13901 2707
rect -13867 2673 -13833 2707
rect -13799 2673 -13765 2707
rect -13731 2673 -13697 2707
rect -13663 2673 -13629 2707
rect -13595 2673 -13561 2707
rect -13527 2673 -13493 2707
rect -13459 2673 -13425 2707
rect -13391 2673 -13357 2707
rect -13323 2673 -13289 2707
rect -13255 2673 -13221 2707
rect -13187 2673 -13153 2707
rect -13119 2673 -13085 2707
rect -13051 2673 -13017 2707
rect -12983 2673 -12949 2707
rect -12915 2673 -12881 2707
rect -12847 2673 -12813 2707
rect -12779 2673 -12745 2707
rect -12711 2673 -12677 2707
rect -12643 2673 -12609 2707
rect -12575 2673 -12541 2707
rect -12507 2673 -12473 2707
rect -12439 2673 -12405 2707
rect -12371 2673 -12337 2707
rect -12303 2673 -12269 2707
rect -12235 2673 -12201 2707
rect -12167 2673 -12133 2707
rect -12099 2673 -12065 2707
rect -12031 2673 -11997 2707
rect -11963 2673 -11929 2707
rect -11895 2673 -11861 2707
rect -11827 2673 -11793 2707
rect -11759 2673 -11725 2707
rect -11691 2673 -11657 2707
rect -11623 2673 -11589 2707
rect -11555 2673 -11521 2707
rect -11487 2673 -11453 2707
rect -11419 2673 -11385 2707
rect -11351 2673 -11317 2707
rect -11283 2673 -11249 2707
rect -11215 2673 -11181 2707
rect -11147 2673 -11113 2707
rect -11079 2673 -11045 2707
rect -11011 2673 -10977 2707
rect -10943 2673 -10909 2707
rect -10875 2673 -10841 2707
rect -10807 2673 -10773 2707
rect -10739 2673 -10705 2707
rect -10671 2673 -10637 2707
rect -10603 2673 -10569 2707
rect -10535 2673 -10501 2707
rect -10467 2673 -10433 2707
rect -10399 2673 -10365 2707
rect -10331 2673 -10297 2707
rect -10263 2673 -10229 2707
rect -10195 2673 -10161 2707
rect -10127 2673 -10093 2707
rect -10059 2673 -10025 2707
rect -9991 2673 -9957 2707
rect -9923 2673 -9889 2707
rect -9855 2673 -9821 2707
rect -9787 2673 -9753 2707
rect -9719 2673 -9685 2707
rect -9651 2673 -9617 2707
rect -9583 2673 -9549 2707
rect -9515 2673 -9481 2707
rect -9447 2673 -9413 2707
<< locali >>
rect -14679 5417 -14521 5451
rect -14487 5417 -14453 5451
rect -14419 5417 -14385 5451
rect -14351 5417 -14317 5451
rect -14283 5417 -14249 5451
rect -14215 5417 -14181 5451
rect -14147 5417 -14113 5451
rect -14079 5417 -14045 5451
rect -14011 5417 -13977 5451
rect -13943 5417 -13909 5451
rect -13875 5417 -13841 5451
rect -13807 5417 -13773 5451
rect -13739 5417 -13705 5451
rect -13671 5417 -13637 5451
rect -13603 5417 -13569 5451
rect -13535 5417 -13501 5451
rect -13467 5417 -13433 5451
rect -13399 5417 -13365 5451
rect -13331 5417 -13297 5451
rect -13263 5417 -13229 5451
rect -13195 5417 -13161 5451
rect -13127 5417 -13093 5451
rect -13059 5417 -13025 5451
rect -12991 5417 -12957 5451
rect -12923 5417 -12889 5451
rect -12855 5417 -12821 5451
rect -12787 5417 -12753 5451
rect -12719 5417 -12685 5451
rect -12651 5417 -12617 5451
rect -12583 5417 -12549 5451
rect -12515 5417 -12481 5451
rect -12447 5417 -12413 5451
rect -12379 5417 -12345 5451
rect -12311 5417 -12277 5451
rect -12243 5417 -12209 5451
rect -12175 5417 -12141 5451
rect -12107 5417 -12073 5451
rect -12039 5417 -12005 5451
rect -11971 5417 -11937 5451
rect -11903 5417 -11869 5451
rect -11835 5417 -11801 5451
rect -11767 5417 -11733 5451
rect -11699 5417 -11665 5451
rect -11631 5417 -11597 5451
rect -11563 5417 -11529 5451
rect -11495 5417 -11461 5451
rect -11427 5417 -11393 5451
rect -11359 5417 -11325 5451
rect -11291 5417 -11257 5451
rect -11223 5417 -11189 5451
rect -11155 5417 -11121 5451
rect -11087 5417 -11053 5451
rect -11019 5417 -10985 5451
rect -10951 5417 -10917 5451
rect -10883 5417 -10849 5451
rect -10815 5417 -10781 5451
rect -10747 5417 -10713 5451
rect -10679 5417 -10645 5451
rect -10611 5417 -10577 5451
rect -10543 5417 -10509 5451
rect -10475 5417 -10441 5451
rect -10407 5417 -10373 5451
rect -10339 5417 -10305 5451
rect -10271 5417 -10237 5451
rect -10203 5417 -10169 5451
rect -10135 5417 -10101 5451
rect -10067 5417 -10033 5451
rect -9999 5417 -9965 5451
rect -9931 5417 -9897 5451
rect -9863 5417 -9829 5451
rect -9795 5417 -9761 5451
rect -9727 5417 -9693 5451
rect -9659 5417 -9625 5451
rect -9591 5417 -9557 5451
rect -9523 5417 -9489 5451
rect -9455 5417 -9193 5451
rect -14679 5251 -14645 5417
rect -14679 5183 -14645 5217
rect -14679 5115 -14645 5149
rect -14679 5047 -14645 5081
rect -14679 4979 -14645 5013
rect -14679 4911 -14645 4945
rect -14679 4843 -14645 4877
rect -14679 4775 -14645 4809
rect -14679 4707 -14645 4741
rect -14679 4639 -14645 4673
rect -14679 4571 -14645 4605
rect -14679 4503 -14645 4537
rect -14679 4435 -14645 4469
rect -14679 4367 -14645 4401
rect -14679 4299 -14645 4333
rect -14679 4231 -14645 4265
rect -14679 4163 -14645 4197
rect -14679 4095 -14645 4129
rect -14679 4027 -14645 4061
rect -14679 3959 -14645 3993
rect -14679 3891 -14645 3925
rect -14679 3823 -14645 3857
rect -14679 3755 -14645 3789
rect -14679 3687 -14645 3721
rect -14679 3619 -14645 3653
rect -14679 3551 -14645 3585
rect -14679 3483 -14645 3517
rect -14679 3415 -14645 3449
rect -14679 3347 -14645 3381
rect -14679 3279 -14645 3313
rect -14679 3211 -14645 3245
rect -14679 3143 -14645 3177
rect -14679 3075 -14645 3109
rect -14679 3007 -14645 3041
rect -14679 2939 -14645 2973
rect -14679 2707 -14645 2905
rect -9227 5251 -9193 5417
rect -9227 5183 -9193 5217
rect -9227 5115 -9193 5149
rect -9227 5047 -9193 5081
rect -9227 4979 -9193 5013
rect -9227 4911 -9193 4945
rect -9227 4843 -9193 4877
rect -9227 4775 -9193 4809
rect -9227 4707 -9193 4741
rect -9227 4639 -9193 4673
rect -9227 4571 -9193 4605
rect -9227 4503 -9193 4537
rect -9227 4435 -9193 4469
rect -9227 4367 -9193 4401
rect -9227 4299 -9193 4333
rect -9227 4231 -9193 4265
rect -9227 4163 -9193 4197
rect -9227 4095 -9193 4129
rect -9227 4027 -9193 4061
rect -9227 3959 -9193 3993
rect -9227 3891 -9193 3925
rect -9227 3823 -9193 3857
rect -9227 3755 -9193 3789
rect -9227 3687 -9193 3721
rect -9227 3619 -9193 3653
rect -9227 3551 -9193 3585
rect -9227 3483 -9193 3517
rect -9227 3415 -9193 3449
rect -9227 3347 -9193 3381
rect -9227 3279 -9193 3313
rect -9227 3211 -9193 3245
rect -9227 3143 -9193 3177
rect -9227 3075 -9193 3109
rect -9227 3007 -9193 3041
rect -9227 2939 -9193 2973
rect -9227 2707 -9193 2905
rect -14679 2673 -14479 2707
rect -14445 2673 -14411 2707
rect -14377 2673 -14343 2707
rect -14309 2673 -14275 2707
rect -14241 2673 -14207 2707
rect -14173 2673 -14139 2707
rect -14105 2673 -14071 2707
rect -14037 2673 -14003 2707
rect -13969 2673 -13935 2707
rect -13901 2673 -13867 2707
rect -13833 2673 -13799 2707
rect -13765 2673 -13731 2707
rect -13697 2673 -13663 2707
rect -13629 2673 -13595 2707
rect -13561 2673 -13527 2707
rect -13493 2673 -13459 2707
rect -13425 2673 -13391 2707
rect -13357 2673 -13323 2707
rect -13289 2673 -13255 2707
rect -13221 2673 -13187 2707
rect -13153 2673 -13119 2707
rect -13085 2673 -13051 2707
rect -13017 2673 -12983 2707
rect -12949 2673 -12915 2707
rect -12881 2673 -12847 2707
rect -12813 2673 -12779 2707
rect -12745 2673 -12711 2707
rect -12677 2673 -12643 2707
rect -12609 2673 -12575 2707
rect -12541 2673 -12507 2707
rect -12473 2673 -12439 2707
rect -12405 2673 -12371 2707
rect -12337 2673 -12303 2707
rect -12269 2673 -12235 2707
rect -12201 2673 -12167 2707
rect -12133 2673 -12099 2707
rect -12065 2673 -12031 2707
rect -11997 2673 -11963 2707
rect -11929 2673 -11895 2707
rect -11861 2673 -11827 2707
rect -11793 2673 -11759 2707
rect -11725 2673 -11691 2707
rect -11657 2673 -11623 2707
rect -11589 2673 -11555 2707
rect -11521 2673 -11487 2707
rect -11453 2673 -11419 2707
rect -11385 2673 -11351 2707
rect -11317 2673 -11283 2707
rect -11249 2673 -11215 2707
rect -11181 2673 -11147 2707
rect -11113 2673 -11079 2707
rect -11045 2673 -11011 2707
rect -10977 2673 -10943 2707
rect -10909 2673 -10875 2707
rect -10841 2673 -10807 2707
rect -10773 2673 -10739 2707
rect -10705 2673 -10671 2707
rect -10637 2673 -10603 2707
rect -10569 2673 -10535 2707
rect -10501 2673 -10467 2707
rect -10433 2673 -10399 2707
rect -10365 2673 -10331 2707
rect -10297 2673 -10263 2707
rect -10229 2673 -10195 2707
rect -10161 2673 -10127 2707
rect -10093 2673 -10059 2707
rect -10025 2673 -9991 2707
rect -9957 2673 -9923 2707
rect -9889 2673 -9855 2707
rect -9821 2673 -9787 2707
rect -9753 2673 -9719 2707
rect -9685 2673 -9651 2707
rect -9617 2673 -9583 2707
rect -9549 2673 -9515 2707
rect -9481 2673 -9447 2707
rect -9413 2673 -9193 2707
<< properties >>
string path -73.520 27.170 -46.050 27.170 -46.050 13.450 -73.310 13.450 -73.310 27.170 
<< end >>
