magic
tech sky130A
magscale 1 2
timestamp 1715010268
<< nwell >>
rect -296 -284 296 284
<< pmos >>
rect -100 -136 100 64
<< pdiff >>
rect -158 49 -100 64
rect -158 15 -146 49
rect -112 15 -100 49
rect -158 -19 -100 15
rect -158 -53 -146 -19
rect -112 -53 -100 -19
rect -158 -87 -100 -53
rect -158 -121 -146 -87
rect -112 -121 -100 -87
rect -158 -136 -100 -121
rect 100 49 158 64
rect 100 15 112 49
rect 146 15 158 49
rect 100 -19 158 15
rect 100 -53 112 -19
rect 146 -53 158 -19
rect 100 -87 158 -53
rect 100 -121 112 -87
rect 146 -121 158 -87
rect 100 -136 158 -121
<< pdiffc >>
rect -146 15 -112 49
rect -146 -53 -112 -19
rect -146 -121 -112 -87
rect 112 15 146 49
rect 112 -53 146 -19
rect 112 -121 146 -87
<< nsubdiff >>
rect -260 214 -153 248
rect -119 214 -85 248
rect -51 214 -17 248
rect 17 214 51 248
rect 85 214 119 248
rect 153 214 260 248
rect -260 119 -226 214
rect -260 51 -226 85
rect 226 119 260 214
rect -260 -17 -226 17
rect -260 -85 -226 -51
rect -260 -214 -226 -119
rect 226 51 260 85
rect 226 -17 260 17
rect 226 -85 260 -51
rect 226 -214 260 -119
rect -260 -248 -153 -214
rect -119 -248 -85 -214
rect -51 -248 -17 -214
rect 17 -248 51 -214
rect 85 -248 119 -214
rect 153 -248 260 -214
<< nsubdiffcont >>
rect -153 214 -119 248
rect -85 214 -51 248
rect -17 214 17 248
rect 51 214 85 248
rect 119 214 153 248
rect -260 85 -226 119
rect 226 85 260 119
rect -260 17 -226 51
rect -260 -51 -226 -17
rect -260 -119 -226 -85
rect 226 17 260 51
rect 226 -51 260 -17
rect 226 -119 260 -85
rect -153 -248 -119 -214
rect -85 -248 -51 -214
rect -17 -248 17 -214
rect 51 -248 85 -214
rect 119 -248 153 -214
<< poly >>
rect -100 145 100 161
rect -100 111 -51 145
rect -17 111 17 145
rect 51 111 100 145
rect -100 64 100 111
rect -100 -162 100 -136
<< polycont >>
rect -51 111 -17 145
rect 17 111 51 145
<< locali >>
rect -260 214 -153 248
rect -119 214 -85 248
rect -51 214 -17 248
rect 17 214 51 248
rect 85 214 119 248
rect 153 214 260 248
rect -260 119 -226 214
rect -100 111 -53 145
rect -17 111 17 145
rect 53 111 100 145
rect 226 119 260 214
rect -260 51 -226 85
rect -260 -17 -226 17
rect -260 -85 -226 -51
rect -260 -214 -226 -119
rect -146 49 -112 68
rect -146 -19 -112 -17
rect -146 -55 -112 -53
rect -146 -140 -112 -121
rect 112 49 146 68
rect 112 -19 146 -17
rect 112 -55 146 -53
rect 112 -140 146 -121
rect 226 51 260 85
rect 226 -17 260 17
rect 226 -85 260 -51
rect 226 -214 260 -119
rect -260 -248 -153 -214
rect -119 -248 -85 -214
rect -51 -248 -17 -214
rect 17 -248 51 -214
rect 85 -248 119 -214
rect 153 -248 260 -214
<< viali >>
rect -53 111 -51 145
rect -51 111 -19 145
rect 19 111 51 145
rect 51 111 53 145
rect -146 15 -112 17
rect -146 -17 -112 15
rect -146 -87 -112 -55
rect -146 -89 -112 -87
rect 112 15 146 17
rect 112 -17 146 15
rect 112 -87 146 -55
rect 112 -89 146 -87
<< metal1 >>
rect -96 145 96 151
rect -96 111 -53 145
rect -19 111 19 145
rect 53 111 96 145
rect -96 105 96 111
rect -152 17 -106 64
rect -152 -17 -146 17
rect -112 -17 -106 17
rect -152 -55 -106 -17
rect -152 -89 -146 -55
rect -112 -89 -106 -55
rect -152 -136 -106 -89
rect 106 17 152 64
rect 106 -17 112 17
rect 146 -17 152 17
rect 106 -55 152 -17
rect 106 -89 112 -55
rect 146 -89 152 -55
rect 106 -136 152 -89
<< properties >>
string FIXED_BBOX -243 -231 243 231
<< end >>
