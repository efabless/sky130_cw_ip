magic
tech sky130A
magscale 1 2
timestamp 1715010268
<< error_p >>
rect -934 5341 48 5403
rect -934 5235 -872 5341
rect -766 5021 -704 5235
rect -766 4959 -120 5021
rect -14 4959 48 5341
<< nwell >>
rect -872 5235 -14 5341
rect -872 4959 -766 5235
rect -120 4959 -14 5235
rect -872 4853 -14 4959
<< nsubdiff >>
rect -836 5271 -749 5305
rect -715 5271 -681 5305
rect -647 5271 -613 5305
rect -579 5271 -545 5305
rect -511 5271 -477 5305
rect -443 5271 -409 5305
rect -375 5271 -341 5305
rect -307 5271 -273 5305
rect -239 5271 -50 5305
rect -836 5165 -802 5271
rect -836 5097 -802 5131
rect -836 4923 -802 5063
rect -84 5165 -50 5271
rect -84 5097 -50 5131
rect -84 4923 -50 5063
rect -836 4889 -696 4923
rect -662 4889 -628 4923
rect -594 4889 -560 4923
rect -526 4889 -492 4923
rect -458 4889 -424 4923
rect -390 4889 -356 4923
rect -322 4889 -288 4923
rect -254 4889 -50 4923
<< nsubdiffcont >>
rect -749 5271 -715 5305
rect -681 5271 -647 5305
rect -613 5271 -579 5305
rect -545 5271 -511 5305
rect -477 5271 -443 5305
rect -409 5271 -375 5305
rect -341 5271 -307 5305
rect -273 5271 -239 5305
rect -836 5131 -802 5165
rect -836 5063 -802 5097
rect -84 5131 -50 5165
rect -84 5063 -50 5097
rect -696 4889 -662 4923
rect -628 4889 -594 4923
rect -560 4889 -526 4923
rect -492 4889 -458 4923
rect -424 4889 -390 4923
rect -356 4889 -322 4923
rect -288 4889 -254 4923
<< locali >>
rect -836 5271 -749 5305
rect -715 5271 -681 5305
rect -647 5271 -613 5305
rect -579 5271 -545 5305
rect -511 5271 -477 5305
rect -443 5271 -409 5305
rect -375 5271 -341 5305
rect -307 5271 -273 5305
rect -239 5271 -50 5305
rect -836 5165 -802 5271
rect -836 5097 -802 5131
rect -836 4923 -802 5063
rect -84 5165 -50 5271
rect -84 5097 -50 5131
rect -84 4923 -50 5063
rect -836 4889 -696 4923
rect -662 4889 -628 4923
rect -594 4889 -560 4923
rect -526 4889 -492 4923
rect -458 4889 -424 4923
rect -390 4889 -356 4923
rect -322 4889 -288 4923
rect -254 4889 -50 4923
<< properties >>
string path -21.800 132.200 -1.675 132.200 -1.675 122.650 -20.475 122.650 -20.475 132.200 
<< end >>
