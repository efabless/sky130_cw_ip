magic
tech sky130A
magscale 1 2
timestamp 1715010268
<< nwell >>
rect 428 -13 13298 3952
<< nsubdiff >>
rect 464 3882 576 3916
rect 610 3882 644 3916
rect 678 3882 712 3916
rect 746 3882 780 3916
rect 814 3882 848 3916
rect 882 3882 916 3916
rect 950 3882 984 3916
rect 1018 3882 1052 3916
rect 1086 3882 1120 3916
rect 1154 3882 1188 3916
rect 1222 3882 1256 3916
rect 1290 3882 1324 3916
rect 1358 3882 1392 3916
rect 1426 3882 1460 3916
rect 1494 3882 1528 3916
rect 1562 3882 1596 3916
rect 1630 3882 1664 3916
rect 1698 3882 1732 3916
rect 1766 3882 1800 3916
rect 1834 3882 1868 3916
rect 1902 3882 1936 3916
rect 1970 3882 2004 3916
rect 2038 3882 2072 3916
rect 2106 3882 2140 3916
rect 2174 3882 2208 3916
rect 2242 3882 2276 3916
rect 2310 3882 2344 3916
rect 2378 3882 2412 3916
rect 2446 3882 2480 3916
rect 2514 3882 2548 3916
rect 2582 3882 2616 3916
rect 2650 3882 2684 3916
rect 2718 3882 2752 3916
rect 2786 3882 2820 3916
rect 2854 3882 2888 3916
rect 2922 3882 2956 3916
rect 2990 3882 3024 3916
rect 3058 3882 3092 3916
rect 3126 3882 3160 3916
rect 3194 3882 3228 3916
rect 3262 3882 3296 3916
rect 3330 3882 3364 3916
rect 3398 3882 3432 3916
rect 3466 3882 3500 3916
rect 3534 3882 3568 3916
rect 3602 3882 3636 3916
rect 3670 3882 3704 3916
rect 3738 3882 3772 3916
rect 3806 3882 3840 3916
rect 3874 3882 3908 3916
rect 3942 3882 3976 3916
rect 4010 3882 4044 3916
rect 4078 3882 4112 3916
rect 4146 3882 4180 3916
rect 4214 3882 4248 3916
rect 4282 3882 4316 3916
rect 4350 3882 4384 3916
rect 4418 3882 4452 3916
rect 4486 3882 4520 3916
rect 4554 3882 4588 3916
rect 4622 3882 4656 3916
rect 4690 3882 4724 3916
rect 4758 3882 4792 3916
rect 4826 3882 4860 3916
rect 4894 3882 4928 3916
rect 4962 3882 4996 3916
rect 5030 3882 5064 3916
rect 5098 3882 5132 3916
rect 5166 3882 5200 3916
rect 5234 3882 5268 3916
rect 5302 3882 5336 3916
rect 5370 3882 5404 3916
rect 5438 3882 5472 3916
rect 5506 3882 5540 3916
rect 5574 3882 5608 3916
rect 5642 3882 5676 3916
rect 5710 3882 5744 3916
rect 5778 3882 5812 3916
rect 5846 3882 5880 3916
rect 5914 3882 5948 3916
rect 5982 3882 6016 3916
rect 6050 3882 6084 3916
rect 6118 3882 6152 3916
rect 6186 3882 6220 3916
rect 6254 3882 6288 3916
rect 6322 3882 6356 3916
rect 6390 3882 6424 3916
rect 6458 3882 6492 3916
rect 6526 3882 6560 3916
rect 6594 3882 6628 3916
rect 6662 3882 6696 3916
rect 6730 3882 6764 3916
rect 6798 3882 6832 3916
rect 6866 3882 6900 3916
rect 6934 3882 6968 3916
rect 7002 3882 7036 3916
rect 7070 3882 7104 3916
rect 7138 3882 7172 3916
rect 7206 3882 7240 3916
rect 7274 3882 7308 3916
rect 7342 3882 7376 3916
rect 7410 3882 7444 3916
rect 7478 3882 7512 3916
rect 7546 3882 7580 3916
rect 7614 3882 7648 3916
rect 7682 3882 7716 3916
rect 7750 3882 7784 3916
rect 7818 3882 7852 3916
rect 7886 3882 7920 3916
rect 7954 3882 7988 3916
rect 8022 3882 8056 3916
rect 8090 3882 8124 3916
rect 8158 3882 8192 3916
rect 8226 3882 8260 3916
rect 8294 3882 8328 3916
rect 8362 3882 8396 3916
rect 8430 3882 8464 3916
rect 8498 3882 8532 3916
rect 8566 3882 8600 3916
rect 8634 3882 8668 3916
rect 8702 3882 8736 3916
rect 8770 3882 8804 3916
rect 8838 3882 8872 3916
rect 8906 3882 8940 3916
rect 8974 3882 9008 3916
rect 9042 3882 9076 3916
rect 9110 3882 9144 3916
rect 9178 3882 9212 3916
rect 9246 3882 9280 3916
rect 9314 3882 9348 3916
rect 9382 3882 9416 3916
rect 9450 3882 9484 3916
rect 9518 3882 9552 3916
rect 9586 3882 9620 3916
rect 9654 3882 9688 3916
rect 9722 3882 9756 3916
rect 9790 3882 9824 3916
rect 9858 3882 9892 3916
rect 9926 3882 9960 3916
rect 9994 3882 10028 3916
rect 10062 3882 10096 3916
rect 10130 3882 10164 3916
rect 10198 3882 10232 3916
rect 10266 3882 10300 3916
rect 10334 3882 10368 3916
rect 10402 3882 10436 3916
rect 10470 3882 10504 3916
rect 10538 3882 10572 3916
rect 10606 3882 10640 3916
rect 10674 3882 10708 3916
rect 10742 3882 10776 3916
rect 10810 3882 10844 3916
rect 10878 3882 10912 3916
rect 10946 3882 10980 3916
rect 11014 3882 11048 3916
rect 11082 3882 11116 3916
rect 11150 3882 11184 3916
rect 11218 3882 11252 3916
rect 11286 3882 11320 3916
rect 11354 3882 11388 3916
rect 11422 3882 11456 3916
rect 11490 3882 11524 3916
rect 11558 3882 11592 3916
rect 11626 3882 11660 3916
rect 11694 3882 11728 3916
rect 11762 3882 11796 3916
rect 11830 3882 11864 3916
rect 11898 3882 11932 3916
rect 11966 3882 12000 3916
rect 12034 3882 12068 3916
rect 12102 3882 12136 3916
rect 12170 3882 12204 3916
rect 12238 3882 12272 3916
rect 12306 3882 12340 3916
rect 12374 3882 12408 3916
rect 12442 3882 12476 3916
rect 12510 3882 12544 3916
rect 12578 3882 12612 3916
rect 12646 3882 12680 3916
rect 12714 3882 12748 3916
rect 12782 3882 12816 3916
rect 12850 3882 12884 3916
rect 12918 3882 12952 3916
rect 12986 3882 13020 3916
rect 13054 3882 13088 3916
rect 13122 3882 13262 3916
rect 464 3776 498 3882
rect 464 3708 498 3742
rect 464 3640 498 3674
rect 464 3572 498 3606
rect 464 3504 498 3538
rect 464 3436 498 3470
rect 464 3368 498 3402
rect 464 3300 498 3334
rect 464 3232 498 3266
rect 464 3164 498 3198
rect 464 3096 498 3130
rect 464 3028 498 3062
rect 464 2960 498 2994
rect 464 2892 498 2926
rect 464 2824 498 2858
rect 464 2756 498 2790
rect 464 2688 498 2722
rect 464 2620 498 2654
rect 464 2552 498 2586
rect 464 2484 498 2518
rect 464 2416 498 2450
rect 464 2348 498 2382
rect 464 2280 498 2314
rect 464 2212 498 2246
rect 464 2144 498 2178
rect 464 2076 498 2110
rect 464 2008 498 2042
rect 464 1940 498 1974
rect 464 1872 498 1906
rect 464 1804 498 1838
rect 464 1736 498 1770
rect 464 1668 498 1702
rect 464 1600 498 1634
rect 464 1532 498 1566
rect 464 1464 498 1498
rect 464 1396 498 1430
rect 464 1328 498 1362
rect 464 1260 498 1294
rect 464 1192 498 1226
rect 464 1124 498 1158
rect 464 1056 498 1090
rect 464 988 498 1022
rect 464 920 498 954
rect 464 852 498 886
rect 464 784 498 818
rect 464 716 498 750
rect 464 648 498 682
rect 464 580 498 614
rect 464 512 498 546
rect 464 444 498 478
rect 464 376 498 410
rect 464 308 498 342
rect 464 240 498 274
rect 464 57 498 206
rect 13228 3776 13262 3882
rect 13228 3708 13262 3742
rect 13228 3640 13262 3674
rect 13228 3572 13262 3606
rect 13228 3504 13262 3538
rect 13228 3436 13262 3470
rect 13228 3368 13262 3402
rect 13228 3300 13262 3334
rect 13228 3232 13262 3266
rect 13228 3164 13262 3198
rect 13228 3096 13262 3130
rect 13228 3028 13262 3062
rect 13228 2960 13262 2994
rect 13228 2892 13262 2926
rect 13228 2824 13262 2858
rect 13228 2756 13262 2790
rect 13228 2688 13262 2722
rect 13228 2620 13262 2654
rect 13228 2552 13262 2586
rect 13228 2484 13262 2518
rect 13228 2416 13262 2450
rect 13228 2348 13262 2382
rect 13228 2280 13262 2314
rect 13228 2212 13262 2246
rect 13228 2144 13262 2178
rect 13228 2076 13262 2110
rect 13228 2008 13262 2042
rect 13228 1940 13262 1974
rect 13228 1872 13262 1906
rect 13228 1804 13262 1838
rect 13228 1736 13262 1770
rect 13228 1668 13262 1702
rect 13228 1600 13262 1634
rect 13228 1532 13262 1566
rect 13228 1464 13262 1498
rect 13228 1396 13262 1430
rect 13228 1328 13262 1362
rect 13228 1260 13262 1294
rect 13228 1192 13262 1226
rect 13228 1124 13262 1158
rect 13228 1056 13262 1090
rect 13228 988 13262 1022
rect 13228 920 13262 954
rect 13228 852 13262 886
rect 13228 784 13262 818
rect 13228 716 13262 750
rect 13228 648 13262 682
rect 13228 580 13262 614
rect 13228 512 13262 546
rect 13228 444 13262 478
rect 13228 376 13262 410
rect 13228 308 13262 342
rect 13228 240 13262 274
rect 13228 57 13262 206
rect 464 23 644 57
rect 678 23 712 57
rect 746 23 780 57
rect 814 23 848 57
rect 882 23 916 57
rect 950 23 984 57
rect 1018 23 1052 57
rect 1086 23 1120 57
rect 1154 23 1188 57
rect 1222 23 1256 57
rect 1290 23 1324 57
rect 1358 23 1392 57
rect 1426 23 1460 57
rect 1494 23 1528 57
rect 1562 23 1596 57
rect 1630 23 1664 57
rect 1698 23 1732 57
rect 1766 23 1800 57
rect 1834 23 1868 57
rect 1902 23 1936 57
rect 1970 23 2004 57
rect 2038 23 2072 57
rect 2106 23 2140 57
rect 2174 23 2208 57
rect 2242 23 2276 57
rect 2310 23 2344 57
rect 2378 23 2412 57
rect 2446 23 2480 57
rect 2514 23 2548 57
rect 2582 23 2616 57
rect 2650 23 2684 57
rect 2718 23 2752 57
rect 2786 23 2820 57
rect 2854 23 2888 57
rect 2922 23 2956 57
rect 2990 23 3024 57
rect 3058 23 3092 57
rect 3126 23 3160 57
rect 3194 23 3228 57
rect 3262 23 3296 57
rect 3330 23 3364 57
rect 3398 23 3432 57
rect 3466 23 3500 57
rect 3534 23 3568 57
rect 3602 23 3636 57
rect 3670 23 3704 57
rect 3738 23 3772 57
rect 3806 23 3840 57
rect 3874 23 3908 57
rect 3942 23 3976 57
rect 4010 23 4044 57
rect 4078 23 4112 57
rect 4146 23 4180 57
rect 4214 23 4248 57
rect 4282 23 4316 57
rect 4350 23 4384 57
rect 4418 23 4452 57
rect 4486 23 4520 57
rect 4554 23 4588 57
rect 4622 23 4656 57
rect 4690 23 4724 57
rect 4758 23 4792 57
rect 4826 23 4860 57
rect 4894 23 4928 57
rect 4962 23 4996 57
rect 5030 23 5064 57
rect 5098 23 5132 57
rect 5166 23 5200 57
rect 5234 23 5268 57
rect 5302 23 5336 57
rect 5370 23 5404 57
rect 5438 23 5472 57
rect 5506 23 5540 57
rect 5574 23 5608 57
rect 5642 23 5676 57
rect 5710 23 5744 57
rect 5778 23 5812 57
rect 5846 23 5880 57
rect 5914 23 5948 57
rect 5982 23 6016 57
rect 6050 23 6084 57
rect 6118 23 6152 57
rect 6186 23 6220 57
rect 6254 23 6288 57
rect 6322 23 6356 57
rect 6390 23 6424 57
rect 6458 23 6492 57
rect 6526 23 6560 57
rect 6594 23 6628 57
rect 6662 23 6696 57
rect 6730 23 6764 57
rect 6798 23 6832 57
rect 6866 23 6900 57
rect 6934 23 6968 57
rect 7002 23 7036 57
rect 7070 23 7104 57
rect 7138 23 7172 57
rect 7206 23 7240 57
rect 7274 23 7308 57
rect 7342 23 7376 57
rect 7410 23 7444 57
rect 7478 23 7512 57
rect 7546 23 7580 57
rect 7614 23 7648 57
rect 7682 23 7716 57
rect 7750 23 7784 57
rect 7818 23 7852 57
rect 7886 23 7920 57
rect 7954 23 7988 57
rect 8022 23 8056 57
rect 8090 23 8124 57
rect 8158 23 8192 57
rect 8226 23 8260 57
rect 8294 23 8328 57
rect 8362 23 8396 57
rect 8430 23 8464 57
rect 8498 23 8532 57
rect 8566 23 8600 57
rect 8634 23 8668 57
rect 8702 23 8736 57
rect 8770 23 8804 57
rect 8838 23 8872 57
rect 8906 23 8940 57
rect 8974 23 9008 57
rect 9042 23 9076 57
rect 9110 23 9144 57
rect 9178 23 9212 57
rect 9246 23 9280 57
rect 9314 23 9348 57
rect 9382 23 9416 57
rect 9450 23 9484 57
rect 9518 23 9552 57
rect 9586 23 9620 57
rect 9654 23 9688 57
rect 9722 23 9756 57
rect 9790 23 9824 57
rect 9858 23 9892 57
rect 9926 23 9960 57
rect 9994 23 10028 57
rect 10062 23 10096 57
rect 10130 23 10164 57
rect 10198 23 10232 57
rect 10266 23 10300 57
rect 10334 23 10368 57
rect 10402 23 10436 57
rect 10470 23 10504 57
rect 10538 23 10572 57
rect 10606 23 10640 57
rect 10674 23 10708 57
rect 10742 23 10776 57
rect 10810 23 10844 57
rect 10878 23 10912 57
rect 10946 23 10980 57
rect 11014 23 11048 57
rect 11082 23 11116 57
rect 11150 23 11184 57
rect 11218 23 11252 57
rect 11286 23 11320 57
rect 11354 23 11388 57
rect 11422 23 11456 57
rect 11490 23 11524 57
rect 11558 23 11592 57
rect 11626 23 11660 57
rect 11694 23 11728 57
rect 11762 23 11796 57
rect 11830 23 11864 57
rect 11898 23 11932 57
rect 11966 23 12000 57
rect 12034 23 12068 57
rect 12102 23 12136 57
rect 12170 23 12204 57
rect 12238 23 12272 57
rect 12306 23 12340 57
rect 12374 23 12408 57
rect 12442 23 12476 57
rect 12510 23 12544 57
rect 12578 23 12612 57
rect 12646 23 12680 57
rect 12714 23 12748 57
rect 12782 23 12816 57
rect 12850 23 12884 57
rect 12918 23 12952 57
rect 12986 23 13020 57
rect 13054 23 13088 57
rect 13122 23 13262 57
<< nsubdiffcont >>
rect 576 3882 610 3916
rect 644 3882 678 3916
rect 712 3882 746 3916
rect 780 3882 814 3916
rect 848 3882 882 3916
rect 916 3882 950 3916
rect 984 3882 1018 3916
rect 1052 3882 1086 3916
rect 1120 3882 1154 3916
rect 1188 3882 1222 3916
rect 1256 3882 1290 3916
rect 1324 3882 1358 3916
rect 1392 3882 1426 3916
rect 1460 3882 1494 3916
rect 1528 3882 1562 3916
rect 1596 3882 1630 3916
rect 1664 3882 1698 3916
rect 1732 3882 1766 3916
rect 1800 3882 1834 3916
rect 1868 3882 1902 3916
rect 1936 3882 1970 3916
rect 2004 3882 2038 3916
rect 2072 3882 2106 3916
rect 2140 3882 2174 3916
rect 2208 3882 2242 3916
rect 2276 3882 2310 3916
rect 2344 3882 2378 3916
rect 2412 3882 2446 3916
rect 2480 3882 2514 3916
rect 2548 3882 2582 3916
rect 2616 3882 2650 3916
rect 2684 3882 2718 3916
rect 2752 3882 2786 3916
rect 2820 3882 2854 3916
rect 2888 3882 2922 3916
rect 2956 3882 2990 3916
rect 3024 3882 3058 3916
rect 3092 3882 3126 3916
rect 3160 3882 3194 3916
rect 3228 3882 3262 3916
rect 3296 3882 3330 3916
rect 3364 3882 3398 3916
rect 3432 3882 3466 3916
rect 3500 3882 3534 3916
rect 3568 3882 3602 3916
rect 3636 3882 3670 3916
rect 3704 3882 3738 3916
rect 3772 3882 3806 3916
rect 3840 3882 3874 3916
rect 3908 3882 3942 3916
rect 3976 3882 4010 3916
rect 4044 3882 4078 3916
rect 4112 3882 4146 3916
rect 4180 3882 4214 3916
rect 4248 3882 4282 3916
rect 4316 3882 4350 3916
rect 4384 3882 4418 3916
rect 4452 3882 4486 3916
rect 4520 3882 4554 3916
rect 4588 3882 4622 3916
rect 4656 3882 4690 3916
rect 4724 3882 4758 3916
rect 4792 3882 4826 3916
rect 4860 3882 4894 3916
rect 4928 3882 4962 3916
rect 4996 3882 5030 3916
rect 5064 3882 5098 3916
rect 5132 3882 5166 3916
rect 5200 3882 5234 3916
rect 5268 3882 5302 3916
rect 5336 3882 5370 3916
rect 5404 3882 5438 3916
rect 5472 3882 5506 3916
rect 5540 3882 5574 3916
rect 5608 3882 5642 3916
rect 5676 3882 5710 3916
rect 5744 3882 5778 3916
rect 5812 3882 5846 3916
rect 5880 3882 5914 3916
rect 5948 3882 5982 3916
rect 6016 3882 6050 3916
rect 6084 3882 6118 3916
rect 6152 3882 6186 3916
rect 6220 3882 6254 3916
rect 6288 3882 6322 3916
rect 6356 3882 6390 3916
rect 6424 3882 6458 3916
rect 6492 3882 6526 3916
rect 6560 3882 6594 3916
rect 6628 3882 6662 3916
rect 6696 3882 6730 3916
rect 6764 3882 6798 3916
rect 6832 3882 6866 3916
rect 6900 3882 6934 3916
rect 6968 3882 7002 3916
rect 7036 3882 7070 3916
rect 7104 3882 7138 3916
rect 7172 3882 7206 3916
rect 7240 3882 7274 3916
rect 7308 3882 7342 3916
rect 7376 3882 7410 3916
rect 7444 3882 7478 3916
rect 7512 3882 7546 3916
rect 7580 3882 7614 3916
rect 7648 3882 7682 3916
rect 7716 3882 7750 3916
rect 7784 3882 7818 3916
rect 7852 3882 7886 3916
rect 7920 3882 7954 3916
rect 7988 3882 8022 3916
rect 8056 3882 8090 3916
rect 8124 3882 8158 3916
rect 8192 3882 8226 3916
rect 8260 3882 8294 3916
rect 8328 3882 8362 3916
rect 8396 3882 8430 3916
rect 8464 3882 8498 3916
rect 8532 3882 8566 3916
rect 8600 3882 8634 3916
rect 8668 3882 8702 3916
rect 8736 3882 8770 3916
rect 8804 3882 8838 3916
rect 8872 3882 8906 3916
rect 8940 3882 8974 3916
rect 9008 3882 9042 3916
rect 9076 3882 9110 3916
rect 9144 3882 9178 3916
rect 9212 3882 9246 3916
rect 9280 3882 9314 3916
rect 9348 3882 9382 3916
rect 9416 3882 9450 3916
rect 9484 3882 9518 3916
rect 9552 3882 9586 3916
rect 9620 3882 9654 3916
rect 9688 3882 9722 3916
rect 9756 3882 9790 3916
rect 9824 3882 9858 3916
rect 9892 3882 9926 3916
rect 9960 3882 9994 3916
rect 10028 3882 10062 3916
rect 10096 3882 10130 3916
rect 10164 3882 10198 3916
rect 10232 3882 10266 3916
rect 10300 3882 10334 3916
rect 10368 3882 10402 3916
rect 10436 3882 10470 3916
rect 10504 3882 10538 3916
rect 10572 3882 10606 3916
rect 10640 3882 10674 3916
rect 10708 3882 10742 3916
rect 10776 3882 10810 3916
rect 10844 3882 10878 3916
rect 10912 3882 10946 3916
rect 10980 3882 11014 3916
rect 11048 3882 11082 3916
rect 11116 3882 11150 3916
rect 11184 3882 11218 3916
rect 11252 3882 11286 3916
rect 11320 3882 11354 3916
rect 11388 3882 11422 3916
rect 11456 3882 11490 3916
rect 11524 3882 11558 3916
rect 11592 3882 11626 3916
rect 11660 3882 11694 3916
rect 11728 3882 11762 3916
rect 11796 3882 11830 3916
rect 11864 3882 11898 3916
rect 11932 3882 11966 3916
rect 12000 3882 12034 3916
rect 12068 3882 12102 3916
rect 12136 3882 12170 3916
rect 12204 3882 12238 3916
rect 12272 3882 12306 3916
rect 12340 3882 12374 3916
rect 12408 3882 12442 3916
rect 12476 3882 12510 3916
rect 12544 3882 12578 3916
rect 12612 3882 12646 3916
rect 12680 3882 12714 3916
rect 12748 3882 12782 3916
rect 12816 3882 12850 3916
rect 12884 3882 12918 3916
rect 12952 3882 12986 3916
rect 13020 3882 13054 3916
rect 13088 3882 13122 3916
rect 464 3742 498 3776
rect 464 3674 498 3708
rect 464 3606 498 3640
rect 464 3538 498 3572
rect 464 3470 498 3504
rect 464 3402 498 3436
rect 464 3334 498 3368
rect 464 3266 498 3300
rect 464 3198 498 3232
rect 464 3130 498 3164
rect 464 3062 498 3096
rect 464 2994 498 3028
rect 464 2926 498 2960
rect 464 2858 498 2892
rect 464 2790 498 2824
rect 464 2722 498 2756
rect 464 2654 498 2688
rect 464 2586 498 2620
rect 464 2518 498 2552
rect 464 2450 498 2484
rect 464 2382 498 2416
rect 464 2314 498 2348
rect 464 2246 498 2280
rect 464 2178 498 2212
rect 464 2110 498 2144
rect 464 2042 498 2076
rect 464 1974 498 2008
rect 464 1906 498 1940
rect 464 1838 498 1872
rect 464 1770 498 1804
rect 464 1702 498 1736
rect 464 1634 498 1668
rect 464 1566 498 1600
rect 464 1498 498 1532
rect 464 1430 498 1464
rect 464 1362 498 1396
rect 464 1294 498 1328
rect 464 1226 498 1260
rect 464 1158 498 1192
rect 464 1090 498 1124
rect 464 1022 498 1056
rect 464 954 498 988
rect 464 886 498 920
rect 464 818 498 852
rect 464 750 498 784
rect 464 682 498 716
rect 464 614 498 648
rect 464 546 498 580
rect 464 478 498 512
rect 464 410 498 444
rect 464 342 498 376
rect 464 274 498 308
rect 464 206 498 240
rect 13228 3742 13262 3776
rect 13228 3674 13262 3708
rect 13228 3606 13262 3640
rect 13228 3538 13262 3572
rect 13228 3470 13262 3504
rect 13228 3402 13262 3436
rect 13228 3334 13262 3368
rect 13228 3266 13262 3300
rect 13228 3198 13262 3232
rect 13228 3130 13262 3164
rect 13228 3062 13262 3096
rect 13228 2994 13262 3028
rect 13228 2926 13262 2960
rect 13228 2858 13262 2892
rect 13228 2790 13262 2824
rect 13228 2722 13262 2756
rect 13228 2654 13262 2688
rect 13228 2586 13262 2620
rect 13228 2518 13262 2552
rect 13228 2450 13262 2484
rect 13228 2382 13262 2416
rect 13228 2314 13262 2348
rect 13228 2246 13262 2280
rect 13228 2178 13262 2212
rect 13228 2110 13262 2144
rect 13228 2042 13262 2076
rect 13228 1974 13262 2008
rect 13228 1906 13262 1940
rect 13228 1838 13262 1872
rect 13228 1770 13262 1804
rect 13228 1702 13262 1736
rect 13228 1634 13262 1668
rect 13228 1566 13262 1600
rect 13228 1498 13262 1532
rect 13228 1430 13262 1464
rect 13228 1362 13262 1396
rect 13228 1294 13262 1328
rect 13228 1226 13262 1260
rect 13228 1158 13262 1192
rect 13228 1090 13262 1124
rect 13228 1022 13262 1056
rect 13228 954 13262 988
rect 13228 886 13262 920
rect 13228 818 13262 852
rect 13228 750 13262 784
rect 13228 682 13262 716
rect 13228 614 13262 648
rect 13228 546 13262 580
rect 13228 478 13262 512
rect 13228 410 13262 444
rect 13228 342 13262 376
rect 13228 274 13262 308
rect 13228 206 13262 240
rect 644 23 678 57
rect 712 23 746 57
rect 780 23 814 57
rect 848 23 882 57
rect 916 23 950 57
rect 984 23 1018 57
rect 1052 23 1086 57
rect 1120 23 1154 57
rect 1188 23 1222 57
rect 1256 23 1290 57
rect 1324 23 1358 57
rect 1392 23 1426 57
rect 1460 23 1494 57
rect 1528 23 1562 57
rect 1596 23 1630 57
rect 1664 23 1698 57
rect 1732 23 1766 57
rect 1800 23 1834 57
rect 1868 23 1902 57
rect 1936 23 1970 57
rect 2004 23 2038 57
rect 2072 23 2106 57
rect 2140 23 2174 57
rect 2208 23 2242 57
rect 2276 23 2310 57
rect 2344 23 2378 57
rect 2412 23 2446 57
rect 2480 23 2514 57
rect 2548 23 2582 57
rect 2616 23 2650 57
rect 2684 23 2718 57
rect 2752 23 2786 57
rect 2820 23 2854 57
rect 2888 23 2922 57
rect 2956 23 2990 57
rect 3024 23 3058 57
rect 3092 23 3126 57
rect 3160 23 3194 57
rect 3228 23 3262 57
rect 3296 23 3330 57
rect 3364 23 3398 57
rect 3432 23 3466 57
rect 3500 23 3534 57
rect 3568 23 3602 57
rect 3636 23 3670 57
rect 3704 23 3738 57
rect 3772 23 3806 57
rect 3840 23 3874 57
rect 3908 23 3942 57
rect 3976 23 4010 57
rect 4044 23 4078 57
rect 4112 23 4146 57
rect 4180 23 4214 57
rect 4248 23 4282 57
rect 4316 23 4350 57
rect 4384 23 4418 57
rect 4452 23 4486 57
rect 4520 23 4554 57
rect 4588 23 4622 57
rect 4656 23 4690 57
rect 4724 23 4758 57
rect 4792 23 4826 57
rect 4860 23 4894 57
rect 4928 23 4962 57
rect 4996 23 5030 57
rect 5064 23 5098 57
rect 5132 23 5166 57
rect 5200 23 5234 57
rect 5268 23 5302 57
rect 5336 23 5370 57
rect 5404 23 5438 57
rect 5472 23 5506 57
rect 5540 23 5574 57
rect 5608 23 5642 57
rect 5676 23 5710 57
rect 5744 23 5778 57
rect 5812 23 5846 57
rect 5880 23 5914 57
rect 5948 23 5982 57
rect 6016 23 6050 57
rect 6084 23 6118 57
rect 6152 23 6186 57
rect 6220 23 6254 57
rect 6288 23 6322 57
rect 6356 23 6390 57
rect 6424 23 6458 57
rect 6492 23 6526 57
rect 6560 23 6594 57
rect 6628 23 6662 57
rect 6696 23 6730 57
rect 6764 23 6798 57
rect 6832 23 6866 57
rect 6900 23 6934 57
rect 6968 23 7002 57
rect 7036 23 7070 57
rect 7104 23 7138 57
rect 7172 23 7206 57
rect 7240 23 7274 57
rect 7308 23 7342 57
rect 7376 23 7410 57
rect 7444 23 7478 57
rect 7512 23 7546 57
rect 7580 23 7614 57
rect 7648 23 7682 57
rect 7716 23 7750 57
rect 7784 23 7818 57
rect 7852 23 7886 57
rect 7920 23 7954 57
rect 7988 23 8022 57
rect 8056 23 8090 57
rect 8124 23 8158 57
rect 8192 23 8226 57
rect 8260 23 8294 57
rect 8328 23 8362 57
rect 8396 23 8430 57
rect 8464 23 8498 57
rect 8532 23 8566 57
rect 8600 23 8634 57
rect 8668 23 8702 57
rect 8736 23 8770 57
rect 8804 23 8838 57
rect 8872 23 8906 57
rect 8940 23 8974 57
rect 9008 23 9042 57
rect 9076 23 9110 57
rect 9144 23 9178 57
rect 9212 23 9246 57
rect 9280 23 9314 57
rect 9348 23 9382 57
rect 9416 23 9450 57
rect 9484 23 9518 57
rect 9552 23 9586 57
rect 9620 23 9654 57
rect 9688 23 9722 57
rect 9756 23 9790 57
rect 9824 23 9858 57
rect 9892 23 9926 57
rect 9960 23 9994 57
rect 10028 23 10062 57
rect 10096 23 10130 57
rect 10164 23 10198 57
rect 10232 23 10266 57
rect 10300 23 10334 57
rect 10368 23 10402 57
rect 10436 23 10470 57
rect 10504 23 10538 57
rect 10572 23 10606 57
rect 10640 23 10674 57
rect 10708 23 10742 57
rect 10776 23 10810 57
rect 10844 23 10878 57
rect 10912 23 10946 57
rect 10980 23 11014 57
rect 11048 23 11082 57
rect 11116 23 11150 57
rect 11184 23 11218 57
rect 11252 23 11286 57
rect 11320 23 11354 57
rect 11388 23 11422 57
rect 11456 23 11490 57
rect 11524 23 11558 57
rect 11592 23 11626 57
rect 11660 23 11694 57
rect 11728 23 11762 57
rect 11796 23 11830 57
rect 11864 23 11898 57
rect 11932 23 11966 57
rect 12000 23 12034 57
rect 12068 23 12102 57
rect 12136 23 12170 57
rect 12204 23 12238 57
rect 12272 23 12306 57
rect 12340 23 12374 57
rect 12408 23 12442 57
rect 12476 23 12510 57
rect 12544 23 12578 57
rect 12612 23 12646 57
rect 12680 23 12714 57
rect 12748 23 12782 57
rect 12816 23 12850 57
rect 12884 23 12918 57
rect 12952 23 12986 57
rect 13020 23 13054 57
rect 13088 23 13122 57
<< locali >>
rect 464 3882 576 3916
rect 610 3882 644 3916
rect 678 3882 712 3916
rect 746 3882 780 3916
rect 814 3882 848 3916
rect 882 3882 916 3916
rect 950 3882 984 3916
rect 1018 3882 1052 3916
rect 1086 3882 1120 3916
rect 1154 3882 1188 3916
rect 1222 3882 1256 3916
rect 1290 3882 1324 3916
rect 1358 3882 1392 3916
rect 1426 3882 1460 3916
rect 1494 3882 1528 3916
rect 1562 3882 1596 3916
rect 1630 3882 1664 3916
rect 1698 3882 1732 3916
rect 1766 3882 1800 3916
rect 1834 3882 1868 3916
rect 1902 3882 1936 3916
rect 1970 3882 2004 3916
rect 2038 3882 2072 3916
rect 2106 3882 2140 3916
rect 2174 3882 2208 3916
rect 2242 3882 2276 3916
rect 2310 3882 2344 3916
rect 2378 3882 2412 3916
rect 2446 3882 2480 3916
rect 2514 3882 2548 3916
rect 2582 3882 2616 3916
rect 2650 3882 2684 3916
rect 2718 3882 2752 3916
rect 2786 3882 2820 3916
rect 2854 3882 2888 3916
rect 2922 3882 2956 3916
rect 2990 3882 3024 3916
rect 3058 3882 3092 3916
rect 3126 3882 3160 3916
rect 3194 3882 3228 3916
rect 3262 3882 3296 3916
rect 3330 3882 3364 3916
rect 3398 3882 3432 3916
rect 3466 3882 3500 3916
rect 3534 3882 3568 3916
rect 3602 3882 3636 3916
rect 3670 3882 3704 3916
rect 3738 3882 3772 3916
rect 3806 3882 3840 3916
rect 3874 3882 3908 3916
rect 3942 3882 3976 3916
rect 4010 3882 4044 3916
rect 4078 3882 4112 3916
rect 4146 3882 4180 3916
rect 4214 3882 4248 3916
rect 4282 3882 4316 3916
rect 4350 3882 4384 3916
rect 4418 3882 4452 3916
rect 4486 3882 4520 3916
rect 4554 3882 4588 3916
rect 4622 3882 4656 3916
rect 4690 3882 4724 3916
rect 4758 3882 4792 3916
rect 4826 3882 4860 3916
rect 4894 3882 4928 3916
rect 4962 3882 4996 3916
rect 5030 3882 5064 3916
rect 5098 3882 5132 3916
rect 5166 3882 5200 3916
rect 5234 3882 5268 3916
rect 5302 3882 5336 3916
rect 5370 3882 5404 3916
rect 5438 3882 5472 3916
rect 5506 3882 5540 3916
rect 5574 3882 5608 3916
rect 5642 3882 5676 3916
rect 5710 3882 5744 3916
rect 5778 3882 5812 3916
rect 5846 3882 5880 3916
rect 5914 3882 5948 3916
rect 5982 3882 6016 3916
rect 6050 3882 6084 3916
rect 6118 3882 6152 3916
rect 6186 3882 6220 3916
rect 6254 3882 6288 3916
rect 6322 3882 6356 3916
rect 6390 3882 6424 3916
rect 6458 3882 6492 3916
rect 6526 3882 6560 3916
rect 6594 3882 6628 3916
rect 6662 3882 6696 3916
rect 6730 3882 6764 3916
rect 6798 3882 6832 3916
rect 6866 3882 6900 3916
rect 6934 3882 6968 3916
rect 7002 3882 7036 3916
rect 7070 3882 7104 3916
rect 7138 3882 7172 3916
rect 7206 3882 7240 3916
rect 7274 3882 7308 3916
rect 7342 3882 7376 3916
rect 7410 3882 7444 3916
rect 7478 3882 7512 3916
rect 7546 3882 7580 3916
rect 7614 3882 7648 3916
rect 7682 3882 7716 3916
rect 7750 3882 7784 3916
rect 7818 3882 7852 3916
rect 7886 3882 7920 3916
rect 7954 3882 7988 3916
rect 8022 3882 8056 3916
rect 8090 3882 8124 3916
rect 8158 3882 8192 3916
rect 8226 3882 8260 3916
rect 8294 3882 8328 3916
rect 8362 3882 8396 3916
rect 8430 3882 8464 3916
rect 8498 3882 8532 3916
rect 8566 3882 8600 3916
rect 8634 3882 8668 3916
rect 8702 3882 8736 3916
rect 8770 3882 8804 3916
rect 8838 3882 8872 3916
rect 8906 3882 8940 3916
rect 8974 3882 9008 3916
rect 9042 3882 9076 3916
rect 9110 3882 9144 3916
rect 9178 3882 9212 3916
rect 9246 3882 9280 3916
rect 9314 3882 9348 3916
rect 9382 3882 9416 3916
rect 9450 3882 9484 3916
rect 9518 3882 9552 3916
rect 9586 3882 9620 3916
rect 9654 3882 9688 3916
rect 9722 3882 9756 3916
rect 9790 3882 9824 3916
rect 9858 3882 9892 3916
rect 9926 3882 9960 3916
rect 9994 3882 10028 3916
rect 10062 3882 10096 3916
rect 10130 3882 10164 3916
rect 10198 3882 10232 3916
rect 10266 3882 10300 3916
rect 10334 3882 10368 3916
rect 10402 3882 10436 3916
rect 10470 3882 10504 3916
rect 10538 3882 10572 3916
rect 10606 3882 10640 3916
rect 10674 3882 10708 3916
rect 10742 3882 10776 3916
rect 10810 3882 10844 3916
rect 10878 3882 10912 3916
rect 10946 3882 10980 3916
rect 11014 3882 11048 3916
rect 11082 3882 11116 3916
rect 11150 3882 11184 3916
rect 11218 3882 11252 3916
rect 11286 3882 11320 3916
rect 11354 3882 11388 3916
rect 11422 3882 11456 3916
rect 11490 3882 11524 3916
rect 11558 3882 11592 3916
rect 11626 3882 11660 3916
rect 11694 3882 11728 3916
rect 11762 3882 11796 3916
rect 11830 3882 11864 3916
rect 11898 3882 11932 3916
rect 11966 3882 12000 3916
rect 12034 3882 12068 3916
rect 12102 3882 12136 3916
rect 12170 3882 12204 3916
rect 12238 3882 12272 3916
rect 12306 3882 12340 3916
rect 12374 3882 12408 3916
rect 12442 3882 12476 3916
rect 12510 3882 12544 3916
rect 12578 3882 12612 3916
rect 12646 3882 12680 3916
rect 12714 3882 12748 3916
rect 12782 3882 12816 3916
rect 12850 3882 12884 3916
rect 12918 3882 12952 3916
rect 12986 3882 13020 3916
rect 13054 3882 13088 3916
rect 13122 3882 13262 3916
rect 464 3776 498 3882
rect 464 3708 498 3742
rect 464 3640 498 3674
rect 464 3572 498 3606
rect 464 3504 498 3538
rect 464 3436 498 3470
rect 464 3368 498 3402
rect 464 3300 498 3334
rect 464 3232 498 3266
rect 464 3164 498 3198
rect 464 3096 498 3130
rect 464 3028 498 3062
rect 464 2960 498 2994
rect 464 2892 498 2926
rect 464 2824 498 2858
rect 464 2756 498 2790
rect 464 2688 498 2722
rect 464 2620 498 2654
rect 464 2552 498 2586
rect 464 2484 498 2518
rect 464 2416 498 2450
rect 464 2348 498 2382
rect 464 2280 498 2314
rect 464 2212 498 2246
rect 464 2144 498 2178
rect 464 2076 498 2110
rect 464 2008 498 2042
rect 464 1940 498 1974
rect 464 1872 498 1906
rect 464 1804 498 1838
rect 464 1736 498 1770
rect 464 1668 498 1702
rect 464 1600 498 1634
rect 464 1532 498 1566
rect 464 1464 498 1498
rect 464 1396 498 1430
rect 464 1328 498 1362
rect 464 1260 498 1294
rect 464 1192 498 1226
rect 464 1124 498 1158
rect 464 1056 498 1090
rect 464 988 498 1022
rect 464 920 498 954
rect 464 852 498 886
rect 464 784 498 818
rect 464 716 498 750
rect 464 648 498 682
rect 464 580 498 614
rect 464 512 498 546
rect 464 444 498 478
rect 464 376 498 410
rect 464 308 498 342
rect 464 240 498 274
rect 464 57 498 206
rect 13228 3776 13262 3882
rect 13228 3708 13262 3742
rect 13228 3640 13262 3674
rect 13228 3572 13262 3606
rect 13228 3504 13262 3538
rect 13228 3436 13262 3470
rect 13228 3368 13262 3402
rect 13228 3300 13262 3334
rect 13228 3232 13262 3266
rect 13228 3164 13262 3198
rect 13228 3096 13262 3130
rect 13228 3028 13262 3062
rect 13228 2960 13262 2994
rect 13228 2892 13262 2926
rect 13228 2824 13262 2858
rect 13228 2756 13262 2790
rect 13228 2688 13262 2722
rect 13228 2620 13262 2654
rect 13228 2552 13262 2586
rect 13228 2484 13262 2518
rect 13228 2416 13262 2450
rect 13228 2348 13262 2382
rect 13228 2280 13262 2314
rect 13228 2212 13262 2246
rect 13228 2144 13262 2178
rect 13228 2076 13262 2110
rect 13228 2008 13262 2042
rect 13228 1940 13262 1974
rect 13228 1872 13262 1906
rect 13228 1804 13262 1838
rect 13228 1736 13262 1770
rect 13228 1668 13262 1702
rect 13228 1600 13262 1634
rect 13228 1532 13262 1566
rect 13228 1464 13262 1498
rect 13228 1396 13262 1430
rect 13228 1328 13262 1362
rect 13228 1260 13262 1294
rect 13228 1192 13262 1226
rect 13228 1124 13262 1158
rect 13228 1056 13262 1090
rect 13228 988 13262 1022
rect 13228 920 13262 954
rect 13228 852 13262 886
rect 13228 784 13262 818
rect 13228 716 13262 750
rect 13228 648 13262 682
rect 13228 580 13262 614
rect 13228 512 13262 546
rect 13228 444 13262 478
rect 13228 376 13262 410
rect 13228 308 13262 342
rect 13228 240 13262 274
rect 13228 57 13262 206
rect 464 23 644 57
rect 678 23 712 57
rect 746 23 780 57
rect 814 23 848 57
rect 882 23 916 57
rect 950 23 984 57
rect 1018 23 1052 57
rect 1086 23 1120 57
rect 1154 23 1188 57
rect 1222 23 1256 57
rect 1290 23 1324 57
rect 1358 23 1392 57
rect 1426 23 1460 57
rect 1494 23 1528 57
rect 1562 23 1596 57
rect 1630 23 1664 57
rect 1698 23 1732 57
rect 1766 23 1800 57
rect 1834 23 1868 57
rect 1902 23 1936 57
rect 1970 23 2004 57
rect 2038 23 2072 57
rect 2106 23 2140 57
rect 2174 23 2208 57
rect 2242 23 2276 57
rect 2310 23 2344 57
rect 2378 23 2412 57
rect 2446 23 2480 57
rect 2514 23 2548 57
rect 2582 23 2616 57
rect 2650 23 2684 57
rect 2718 23 2752 57
rect 2786 23 2820 57
rect 2854 23 2888 57
rect 2922 23 2956 57
rect 2990 23 3024 57
rect 3058 23 3092 57
rect 3126 23 3160 57
rect 3194 23 3228 57
rect 3262 23 3296 57
rect 3330 23 3364 57
rect 3398 23 3432 57
rect 3466 23 3500 57
rect 3534 23 3568 57
rect 3602 23 3636 57
rect 3670 23 3704 57
rect 3738 23 3772 57
rect 3806 23 3840 57
rect 3874 23 3908 57
rect 3942 23 3976 57
rect 4010 23 4044 57
rect 4078 23 4112 57
rect 4146 23 4180 57
rect 4214 23 4248 57
rect 4282 23 4316 57
rect 4350 23 4384 57
rect 4418 23 4452 57
rect 4486 23 4520 57
rect 4554 23 4588 57
rect 4622 23 4656 57
rect 4690 23 4724 57
rect 4758 23 4792 57
rect 4826 23 4860 57
rect 4894 23 4928 57
rect 4962 23 4996 57
rect 5030 23 5064 57
rect 5098 23 5132 57
rect 5166 23 5200 57
rect 5234 23 5268 57
rect 5302 23 5336 57
rect 5370 23 5404 57
rect 5438 23 5472 57
rect 5506 23 5540 57
rect 5574 23 5608 57
rect 5642 23 5676 57
rect 5710 23 5744 57
rect 5778 23 5812 57
rect 5846 23 5880 57
rect 5914 23 5948 57
rect 5982 23 6016 57
rect 6050 23 6084 57
rect 6118 23 6152 57
rect 6186 23 6220 57
rect 6254 23 6288 57
rect 6322 23 6356 57
rect 6390 23 6424 57
rect 6458 23 6492 57
rect 6526 23 6560 57
rect 6594 23 6628 57
rect 6662 23 6696 57
rect 6730 23 6764 57
rect 6798 23 6832 57
rect 6866 23 6900 57
rect 6934 23 6968 57
rect 7002 23 7036 57
rect 7070 23 7104 57
rect 7138 23 7172 57
rect 7206 23 7240 57
rect 7274 23 7308 57
rect 7342 23 7376 57
rect 7410 23 7444 57
rect 7478 23 7512 57
rect 7546 23 7580 57
rect 7614 23 7648 57
rect 7682 23 7716 57
rect 7750 23 7784 57
rect 7818 23 7852 57
rect 7886 23 7920 57
rect 7954 23 7988 57
rect 8022 23 8056 57
rect 8090 23 8124 57
rect 8158 23 8192 57
rect 8226 23 8260 57
rect 8294 23 8328 57
rect 8362 23 8396 57
rect 8430 23 8464 57
rect 8498 23 8532 57
rect 8566 23 8600 57
rect 8634 23 8668 57
rect 8702 23 8736 57
rect 8770 23 8804 57
rect 8838 23 8872 57
rect 8906 23 8940 57
rect 8974 23 9008 57
rect 9042 23 9076 57
rect 9110 23 9144 57
rect 9178 23 9212 57
rect 9246 23 9280 57
rect 9314 23 9348 57
rect 9382 23 9416 57
rect 9450 23 9484 57
rect 9518 23 9552 57
rect 9586 23 9620 57
rect 9654 23 9688 57
rect 9722 23 9756 57
rect 9790 23 9824 57
rect 9858 23 9892 57
rect 9926 23 9960 57
rect 9994 23 10028 57
rect 10062 23 10096 57
rect 10130 23 10164 57
rect 10198 23 10232 57
rect 10266 23 10300 57
rect 10334 23 10368 57
rect 10402 23 10436 57
rect 10470 23 10504 57
rect 10538 23 10572 57
rect 10606 23 10640 57
rect 10674 23 10708 57
rect 10742 23 10776 57
rect 10810 23 10844 57
rect 10878 23 10912 57
rect 10946 23 10980 57
rect 11014 23 11048 57
rect 11082 23 11116 57
rect 11150 23 11184 57
rect 11218 23 11252 57
rect 11286 23 11320 57
rect 11354 23 11388 57
rect 11422 23 11456 57
rect 11490 23 11524 57
rect 11558 23 11592 57
rect 11626 23 11660 57
rect 11694 23 11728 57
rect 11762 23 11796 57
rect 11830 23 11864 57
rect 11898 23 11932 57
rect 11966 23 12000 57
rect 12034 23 12068 57
rect 12102 23 12136 57
rect 12170 23 12204 57
rect 12238 23 12272 57
rect 12306 23 12340 57
rect 12374 23 12408 57
rect 12442 23 12476 57
rect 12510 23 12544 57
rect 12578 23 12612 57
rect 12646 23 12680 57
rect 12714 23 12748 57
rect 12782 23 12816 57
rect 12850 23 12884 57
rect 12918 23 12952 57
rect 12986 23 13020 57
rect 13054 23 13088 57
rect 13122 23 13262 57
<< properties >>
string path 2.140 19.495 66.225 19.495 66.225 0.200 2.405 0.200 2.405 19.495 
<< end >>
