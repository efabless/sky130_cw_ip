magic
tech sky130A
magscale 1 2
timestamp 1715010268
<< pwell >>
rect -236 -369 236 369
<< nmos >>
rect -50 -231 50 169
<< ndiff >>
rect -108 156 -50 169
rect -108 122 -96 156
rect -62 122 -50 156
rect -108 88 -50 122
rect -108 54 -96 88
rect -62 54 -50 88
rect -108 20 -50 54
rect -108 -14 -96 20
rect -62 -14 -50 20
rect -108 -48 -50 -14
rect -108 -82 -96 -48
rect -62 -82 -50 -48
rect -108 -116 -50 -82
rect -108 -150 -96 -116
rect -62 -150 -50 -116
rect -108 -184 -50 -150
rect -108 -218 -96 -184
rect -62 -218 -50 -184
rect -108 -231 -50 -218
rect 50 156 108 169
rect 50 122 62 156
rect 96 122 108 156
rect 50 88 108 122
rect 50 54 62 88
rect 96 54 108 88
rect 50 20 108 54
rect 50 -14 62 20
rect 96 -14 108 20
rect 50 -48 108 -14
rect 50 -82 62 -48
rect 96 -82 108 -48
rect 50 -116 108 -82
rect 50 -150 62 -116
rect 96 -150 108 -116
rect 50 -184 108 -150
rect 50 -218 62 -184
rect 96 -218 108 -184
rect 50 -231 108 -218
<< ndiffc >>
rect -96 122 -62 156
rect -96 54 -62 88
rect -96 -14 -62 20
rect -96 -82 -62 -48
rect -96 -150 -62 -116
rect -96 -218 -62 -184
rect 62 122 96 156
rect 62 54 96 88
rect 62 -14 96 20
rect 62 -82 96 -48
rect 62 -150 96 -116
rect 62 -218 96 -184
<< psubdiff >>
rect -210 309 -85 343
rect -51 309 -17 343
rect 17 309 51 343
rect 85 309 210 343
rect -210 221 -176 309
rect -210 153 -176 187
rect 176 221 210 309
rect -210 85 -176 119
rect -210 17 -176 51
rect -210 -51 -176 -17
rect -210 -119 -176 -85
rect -210 -187 -176 -153
rect -210 -309 -176 -221
rect 176 153 210 187
rect 176 85 210 119
rect 176 17 210 51
rect 176 -51 210 -17
rect 176 -119 210 -85
rect 176 -187 210 -153
rect 176 -309 210 -221
rect -210 -343 -85 -309
rect -51 -343 -17 -309
rect 17 -343 51 -309
rect 85 -343 210 -309
<< psubdiffcont >>
rect -85 309 -51 343
rect -17 309 17 343
rect 51 309 85 343
rect -210 187 -176 221
rect 176 187 210 221
rect -210 119 -176 153
rect -210 51 -176 85
rect -210 -17 -176 17
rect -210 -85 -176 -51
rect -210 -153 -176 -119
rect -210 -221 -176 -187
rect 176 119 210 153
rect 176 51 210 85
rect 176 -17 210 17
rect 176 -85 210 -51
rect 176 -153 210 -119
rect 176 -221 210 -187
rect -85 -343 -51 -309
rect -17 -343 17 -309
rect 51 -343 85 -309
<< poly >>
rect -50 241 50 257
rect -50 207 -17 241
rect 17 207 50 241
rect -50 169 50 207
rect -50 -257 50 -231
<< polycont >>
rect -17 207 17 241
<< locali >>
rect -210 309 -85 343
rect -51 309 -17 343
rect 17 309 51 343
rect 85 309 210 343
rect -210 221 -176 309
rect -50 207 -17 241
rect 17 207 50 241
rect 176 221 210 309
rect -210 153 -176 187
rect -210 85 -176 119
rect -210 17 -176 51
rect -210 -51 -176 -17
rect -210 -119 -176 -85
rect -210 -187 -176 -153
rect -210 -309 -176 -221
rect -96 156 -62 173
rect -96 88 -62 96
rect -96 20 -62 24
rect -96 -86 -62 -82
rect -96 -158 -62 -150
rect -96 -235 -62 -218
rect 62 156 96 173
rect 62 88 96 96
rect 62 20 96 24
rect 62 -86 96 -82
rect 62 -158 96 -150
rect 62 -235 96 -218
rect 176 153 210 187
rect 176 85 210 119
rect 176 17 210 51
rect 176 -51 210 -17
rect 176 -119 210 -85
rect 176 -187 210 -153
rect 176 -309 210 -221
rect -210 -343 -85 -309
rect -51 -343 -17 -309
rect 17 -343 51 -309
rect 85 -343 210 -309
<< viali >>
rect -17 207 17 241
rect -96 122 -62 130
rect -96 96 -62 122
rect -96 54 -62 58
rect -96 24 -62 54
rect -96 -48 -62 -14
rect -96 -116 -62 -86
rect -96 -120 -62 -116
rect -96 -184 -62 -158
rect -96 -192 -62 -184
rect 62 122 96 130
rect 62 96 96 122
rect 62 54 96 58
rect 62 24 96 54
rect 62 -48 96 -14
rect 62 -116 96 -86
rect 62 -120 96 -116
rect 62 -184 96 -158
rect 62 -192 96 -184
<< metal1 >>
rect -46 241 46 247
rect -46 207 -17 241
rect 17 207 46 241
rect -46 201 46 207
rect -102 130 -56 169
rect -102 96 -96 130
rect -62 96 -56 130
rect -102 58 -56 96
rect -102 24 -96 58
rect -62 24 -56 58
rect -102 -14 -56 24
rect -102 -48 -96 -14
rect -62 -48 -56 -14
rect -102 -86 -56 -48
rect -102 -120 -96 -86
rect -62 -120 -56 -86
rect -102 -158 -56 -120
rect -102 -192 -96 -158
rect -62 -192 -56 -158
rect -102 -231 -56 -192
rect 56 130 102 169
rect 56 96 62 130
rect 96 96 102 130
rect 56 58 102 96
rect 56 24 62 58
rect 96 24 102 58
rect 56 -14 102 24
rect 56 -48 62 -14
rect 96 -48 102 -14
rect 56 -86 102 -48
rect 56 -120 62 -86
rect 96 -120 102 -86
rect 56 -158 102 -120
rect 56 -192 62 -158
rect 96 -192 102 -158
rect 56 -231 102 -192
<< properties >>
string FIXED_BBOX -193 -326 193 326
<< end >>
