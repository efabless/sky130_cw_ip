magic
tech sky130A
magscale 1 2
timestamp 1715010268
<< pwell >>
rect 1438 1395 4377 1481
rect 1438 719 1524 1395
rect 4291 719 4377 1395
rect 1438 633 4377 719
<< psubdiff >>
rect 1464 1421 1669 1455
rect 1703 1421 1737 1455
rect 1771 1421 1805 1455
rect 1839 1421 1873 1455
rect 1907 1421 1941 1455
rect 1975 1421 2009 1455
rect 2043 1421 2077 1455
rect 2111 1421 2145 1455
rect 2179 1421 2213 1455
rect 2247 1421 2281 1455
rect 2315 1421 2349 1455
rect 2383 1421 2417 1455
rect 2451 1421 2485 1455
rect 2519 1421 2553 1455
rect 2587 1421 2621 1455
rect 2655 1421 2689 1455
rect 2723 1421 2757 1455
rect 2791 1421 2825 1455
rect 2859 1421 2893 1455
rect 2927 1421 2961 1455
rect 2995 1421 3029 1455
rect 3063 1421 3097 1455
rect 3131 1421 3165 1455
rect 3199 1421 3233 1455
rect 3267 1421 3301 1455
rect 3335 1421 3369 1455
rect 3403 1421 3437 1455
rect 3471 1421 3505 1455
rect 3539 1421 3573 1455
rect 3607 1421 3641 1455
rect 3675 1421 3709 1455
rect 3743 1421 3777 1455
rect 3811 1421 3845 1455
rect 3879 1421 3913 1455
rect 3947 1421 3981 1455
rect 4015 1421 4049 1455
rect 4083 1421 4117 1455
rect 4151 1421 4351 1455
rect 1464 1255 1498 1421
rect 1464 1187 1498 1221
rect 1464 1119 1498 1153
rect 1464 1051 1498 1085
rect 1464 983 1498 1017
rect 1464 915 1498 949
rect 1464 693 1498 881
rect 4317 1255 4351 1421
rect 4317 1187 4351 1221
rect 4317 1119 4351 1153
rect 4317 1051 4351 1085
rect 4317 983 4351 1017
rect 4317 915 4351 949
rect 4317 693 4351 881
rect 1464 659 1669 693
rect 1703 659 1737 693
rect 1771 659 1805 693
rect 1839 659 1873 693
rect 1907 659 1941 693
rect 1975 659 2009 693
rect 2043 659 2077 693
rect 2111 659 2145 693
rect 2179 659 2213 693
rect 2247 659 2281 693
rect 2315 659 2349 693
rect 2383 659 2417 693
rect 2451 659 2485 693
rect 2519 659 2553 693
rect 2587 659 2621 693
rect 2655 659 2689 693
rect 2723 659 2757 693
rect 2791 659 2825 693
rect 2859 659 2893 693
rect 2927 659 2961 693
rect 2995 659 3029 693
rect 3063 659 3097 693
rect 3131 659 3165 693
rect 3199 659 3233 693
rect 3267 659 3301 693
rect 3335 659 3369 693
rect 3403 659 3437 693
rect 3471 659 3505 693
rect 3539 659 3573 693
rect 3607 659 3641 693
rect 3675 659 3709 693
rect 3743 659 3777 693
rect 3811 659 3845 693
rect 3879 659 3913 693
rect 3947 659 3981 693
rect 4015 659 4049 693
rect 4083 659 4117 693
rect 4151 659 4351 693
<< psubdiffcont >>
rect 1669 1421 1703 1455
rect 1737 1421 1771 1455
rect 1805 1421 1839 1455
rect 1873 1421 1907 1455
rect 1941 1421 1975 1455
rect 2009 1421 2043 1455
rect 2077 1421 2111 1455
rect 2145 1421 2179 1455
rect 2213 1421 2247 1455
rect 2281 1421 2315 1455
rect 2349 1421 2383 1455
rect 2417 1421 2451 1455
rect 2485 1421 2519 1455
rect 2553 1421 2587 1455
rect 2621 1421 2655 1455
rect 2689 1421 2723 1455
rect 2757 1421 2791 1455
rect 2825 1421 2859 1455
rect 2893 1421 2927 1455
rect 2961 1421 2995 1455
rect 3029 1421 3063 1455
rect 3097 1421 3131 1455
rect 3165 1421 3199 1455
rect 3233 1421 3267 1455
rect 3301 1421 3335 1455
rect 3369 1421 3403 1455
rect 3437 1421 3471 1455
rect 3505 1421 3539 1455
rect 3573 1421 3607 1455
rect 3641 1421 3675 1455
rect 3709 1421 3743 1455
rect 3777 1421 3811 1455
rect 3845 1421 3879 1455
rect 3913 1421 3947 1455
rect 3981 1421 4015 1455
rect 4049 1421 4083 1455
rect 4117 1421 4151 1455
rect 1464 1221 1498 1255
rect 1464 1153 1498 1187
rect 1464 1085 1498 1119
rect 1464 1017 1498 1051
rect 1464 949 1498 983
rect 1464 881 1498 915
rect 4317 1221 4351 1255
rect 4317 1153 4351 1187
rect 4317 1085 4351 1119
rect 4317 1017 4351 1051
rect 4317 949 4351 983
rect 4317 881 4351 915
rect 1669 659 1703 693
rect 1737 659 1771 693
rect 1805 659 1839 693
rect 1873 659 1907 693
rect 1941 659 1975 693
rect 2009 659 2043 693
rect 2077 659 2111 693
rect 2145 659 2179 693
rect 2213 659 2247 693
rect 2281 659 2315 693
rect 2349 659 2383 693
rect 2417 659 2451 693
rect 2485 659 2519 693
rect 2553 659 2587 693
rect 2621 659 2655 693
rect 2689 659 2723 693
rect 2757 659 2791 693
rect 2825 659 2859 693
rect 2893 659 2927 693
rect 2961 659 2995 693
rect 3029 659 3063 693
rect 3097 659 3131 693
rect 3165 659 3199 693
rect 3233 659 3267 693
rect 3301 659 3335 693
rect 3369 659 3403 693
rect 3437 659 3471 693
rect 3505 659 3539 693
rect 3573 659 3607 693
rect 3641 659 3675 693
rect 3709 659 3743 693
rect 3777 659 3811 693
rect 3845 659 3879 693
rect 3913 659 3947 693
rect 3981 659 4015 693
rect 4049 659 4083 693
rect 4117 659 4151 693
<< locali >>
rect 1464 1421 1669 1455
rect 1703 1421 1737 1455
rect 1771 1421 1805 1455
rect 1839 1421 1873 1455
rect 1907 1421 1941 1455
rect 1975 1421 2009 1455
rect 2043 1421 2077 1455
rect 2111 1421 2145 1455
rect 2179 1421 2213 1455
rect 2247 1421 2281 1455
rect 2315 1421 2349 1455
rect 2383 1421 2417 1455
rect 2451 1421 2485 1455
rect 2519 1421 2553 1455
rect 2587 1421 2621 1455
rect 2655 1421 2689 1455
rect 2723 1421 2757 1455
rect 2791 1421 2825 1455
rect 2859 1421 2893 1455
rect 2927 1421 2961 1455
rect 2995 1421 3029 1455
rect 3063 1421 3097 1455
rect 3131 1421 3165 1455
rect 3199 1421 3233 1455
rect 3267 1421 3301 1455
rect 3335 1421 3369 1455
rect 3403 1421 3437 1455
rect 3471 1421 3505 1455
rect 3539 1421 3573 1455
rect 3607 1421 3641 1455
rect 3675 1421 3709 1455
rect 3743 1421 3777 1455
rect 3811 1421 3845 1455
rect 3879 1421 3913 1455
rect 3947 1421 3981 1455
rect 4015 1421 4049 1455
rect 4083 1421 4117 1455
rect 4151 1421 4351 1455
rect 1464 1255 1498 1421
rect 1464 1187 1498 1221
rect 1464 1119 1498 1153
rect 1464 1051 1498 1085
rect 1464 983 1498 1017
rect 1464 915 1498 949
rect 1464 693 1498 881
rect 4317 1255 4351 1421
rect 4317 1187 4351 1221
rect 4317 1119 4351 1153
rect 4317 1051 4351 1085
rect 4317 983 4351 1017
rect 4317 915 4351 949
rect 4317 693 4351 881
rect 1464 659 1669 693
rect 1703 659 1737 693
rect 1771 659 1805 693
rect 1839 659 1873 693
rect 1907 659 1941 693
rect 1975 659 2009 693
rect 2043 659 2077 693
rect 2111 659 2145 693
rect 2179 659 2213 693
rect 2247 659 2281 693
rect 2315 659 2349 693
rect 2383 659 2417 693
rect 2451 659 2485 693
rect 2519 659 2553 693
rect 2587 659 2621 693
rect 2655 659 2689 693
rect 2723 659 2757 693
rect 2791 659 2825 693
rect 2859 659 2893 693
rect 2927 659 2961 693
rect 2995 659 3029 693
rect 3063 659 3097 693
rect 3131 659 3165 693
rect 3199 659 3233 693
rect 3267 659 3301 693
rect 3335 659 3369 693
rect 3403 659 3437 693
rect 3471 659 3505 693
rect 3539 659 3573 693
rect 3607 659 3641 693
rect 3675 659 3709 693
rect 3743 659 3777 693
rect 3811 659 3845 693
rect 3879 659 3913 693
rect 3947 659 3981 693
rect 4015 659 4049 693
rect 4083 659 4117 693
rect 4151 659 4351 693
<< properties >>
string path 35.975 35.950 108.350 35.950 108.350 16.900 37.025 16.900 37.025 35.950 
<< end >>
